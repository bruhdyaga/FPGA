`ifndef FACQ_PRN_GEN_SVH
`define FACQ_PRN_GEN_SVH

localparam FACQ_PRNSIZE           = 14;
localparam FACQ_CNTRSIZE          = 23;

localparam FACQ_GPS_L5_PATTERN = 13'b1011111111111;

`endif
