/* `define CRPA_NUMB         2

`define CRPA_HETERODYNE
`define CRPA_UP_HETERODYNE
// `define HETERODYNE_RECORDER
// `define HETERODYNE_DATCOLL
`define HETERODYNE_FIR_ORDER  10

// `define CRPA_DATCOLL

// `define CRPA_D_WIDTH      14
// `define CRPA_C_WIDTH      14
// `define CRPA_ANT          4
// `define CRPA_NCH          (`CRPA_ANT `ifdef CRPA_HETERODYNE * 2 `endif)
// `define CRPA_NT           4
// `define CRPA_NNF          1
`define CRPA_ACCUM_WIDTH  48
`define RAM_SIZE          10  // 2^RAM_SIZE
`define RAM_BLOCKS        40  // numbers from 1 */
