`timescale 1ns / 1ps

module randn_u(
    //.number(0)       // Порядковый номер блока (отличаются зерном)
    // ) insname (
    clk, 
    reset_n, 
    out
    );
    
    parameter number = 0;
    
    input clk;
    input reset_n;
    output out;
    
    wire clk;
    wire reset_n;
    reg [7:0] out;
    
    reg [7:0] X_1;
    reg [7:0] X_2;
    reg [7:0] X_3;
    reg [7:0] X_4;
    reg [7:0] X_5;
    reg [7:0] X_6;
    reg [7:0] X_7;
    reg [7:0] X_8;
    reg [7:0] X_9;
    reg [7:0] X_10;
    reg [7:0] X_11;
    reg [7:0] X_12;
    reg [7:0] X_13;
    reg [7:0] X_14;
    reg [7:0] X_15;
    reg [7:0] X_16;
    reg [7:0] X_17;
    reg [7:0] X_18;
    reg [7:0] X_19;
    reg [7:0] X_20;
    reg [7:0] X_21;
    reg [7:0] X_22;
    reg [7:0] X_23;
    reg [7:0] X_24;
    reg [7:0] X_25;
    reg [7:0] X_26;
    reg [7:0] X_27;
    reg [7:0] X_28;
    reg [7:0] X_29;
    reg [7:0] X_30;
    reg [7:0] X_31;
    reg [7:0] X_32;
    reg [7:0] X_33;
    reg [7:0] X_34;
    reg [7:0] X_35;
    reg [7:0] X_36;
    reg [7:0] X_37;
    reg [7:0] X_38;
    reg [7:0] X_39;
    reg [7:0] X_40;
    reg [7:0] X_41;
    reg [7:0] X_42;
    reg [7:0] X_43;
    reg [7:0] X_44;
    reg [7:0] X_45;
    reg [7:0] X_46;
    reg [7:0] X_47;
    reg [7:0] X_48;
    reg [7:0] X_49;
    reg [7:0] X_50;
    reg [7:0] X_51;
    reg [7:0] X_52;
    reg [7:0] X_53;
    reg [7:0] X_54;
    reg [7:0] X_55;

    always @(posedge clk or negedge reset_n) begin
        if (reset_n == 0) begin
        
            if (number == 0) begin
                X_1 <= 208;
                X_2 <= 231;
                X_3 <= 32;
                X_4 <= 233;
                X_5 <= 161;
                X_6 <= 24;
                X_7 <= 71;
                X_8 <= 140;
                X_9 <= 245;
                X_10 <= 247;
                X_11 <= 40;
                X_12 <= 248;
                X_13 <= 245;
                X_14 <= 124;
                X_15 <= 204;
                X_16 <= 36;
                X_17 <= 107;
                X_18 <= 234;
                X_19 <= 202;
                X_20 <= 245;
                X_21 <= 167;
                X_22 <= 9;
                X_23 <= 217;
                X_24 <= 239;
                X_25 <= 173;
                X_26 <= 193;
                X_27 <= 190;
                X_28 <= 100;
                X_29 <= 167;
                X_30 <= 43;
                X_31 <= 180;
                X_32 <= 8;
                X_33 <= 70;
                X_34 <= 11;
                X_35 <= 24;
                X_36 <= 210;
                X_37 <= 177;
                X_38 <= 81;
                X_39 <= 243;
                X_40 <= 8;
                X_41 <= 112;
                X_42 <= 97;
                X_43 <= 195;
                X_44 <= 203;
                X_45 <= 47;
                X_46 <= 125;
                X_47 <= 114;
                X_48 <= 165;
                X_49 <= 181;
                X_50 <= 193;
                X_51 <= 70;
                X_52 <= 174;
                X_53 <= 167;
                X_54 <= 41;
                X_55 <= 30;
                out <= 0;
            end else if (number == 1) begin
                X_1 <= 127;
                X_2 <= 245;
                X_3 <= 87;
                X_4 <= 149;
                X_5 <= 57;
                X_6 <= 192;
                X_7 <= 65;
                X_8 <= 129;
                X_9 <= 178;
                X_10 <= 228;
                X_11 <= 245;
                X_12 <= 140;
                X_13 <= 35;
                X_14 <= 38;
                X_15 <= 65;
                X_16 <= 215;
                X_17 <= 65;
                X_18 <= 208;
                X_19 <= 62;
                X_20 <= 237;
                X_21 <= 89;
                X_22 <= 50;
                X_23 <= 64;
                X_24 <= 157;
                X_25 <= 121;
                X_26 <= 90;
                X_27 <= 212;
                X_28 <= 149;
                X_29 <= 140;
                X_30 <= 234;
                X_31 <= 73;
                X_32 <= 193;
                X_33 <= 192;
                X_34 <= 97;
                X_35 <= 145;
                X_36 <= 19;
                X_37 <= 13;
                X_38 <= 135;
                X_39 <= 199;
                X_40 <= 239;
                X_41 <= 33;
                X_42 <= 145;
                X_43 <= 120;
                X_44 <= 3;
                X_45 <= 86;
                X_46 <= 41;
                X_47 <= 203;
                X_48 <= 79;
                X_49 <= 135;
                X_50 <= 42;
                X_51 <= 154;
                X_52 <= 67;
                X_53 <= 167;
                X_54 <= 176;
                X_55 <= 191;
                out <= 0;
            end else if (number == 2) begin
                X_1 <= 115;
                X_2 <= 21;
                X_3 <= 58;
                X_4 <= 233;
                X_5 <= 39;
                X_6 <= 211;
                X_7 <= 137;
                X_8 <= 255;
                X_9 <= 20;
                X_10 <= 113;
                X_11 <= 27;
                X_12 <= 246;
                X_13 <= 1;
                X_14 <= 198;
                X_15 <= 209;
                X_16 <= 222;
                X_17 <= 21;
                X_18 <= 102;
                X_19 <= 66;
                X_20 <= 204;
                X_21 <= 110;
                X_22 <= 233;
                X_23 <= 46;
                X_24 <= 67;
                X_25 <= 37;
                X_26 <= 34;
                X_27 <= 222;
                X_28 <= 148;
                X_29 <= 140;
                X_30 <= 37;
                X_31 <= 218;
                X_32 <= 159;
                X_33 <= 89;
                X_34 <= 131;
                X_35 <= 102;
                X_36 <= 19;
                X_37 <= 61;
                X_38 <= 31;
                X_39 <= 47;
                X_40 <= 61;
                X_41 <= 106;
                X_42 <= 12;
                X_43 <= 231;
                X_44 <= 241;
                X_45 <= 125;
                X_46 <= 125;
                X_47 <= 86;
                X_48 <= 230;
                X_49 <= 94;
                X_50 <= 28;
                X_51 <= 199;
                X_52 <= 99;
                X_53 <= 61;
                X_54 <= 103;
                X_55 <= 24;
                out <= 0;
            end else if (number == 3) begin
                X_1 <= 33;
                X_2 <= 241;
                X_3 <= 244;
                X_4 <= 147;
                X_5 <= 15;
                X_6 <= 60;
                X_7 <= 90;
                X_8 <= 210;
                X_9 <= 3;
                X_10 <= 11;
                X_11 <= 43;
                X_12 <= 166;
                X_13 <= 187;
                X_14 <= 165;
                X_15 <= 115;
                X_16 <= 140;
                X_17 <= 75;
                X_18 <= 190;
                X_19 <= 48;
                X_20 <= 175;
                X_21 <= 46;
                X_22 <= 94;
                X_23 <= 160;
                X_24 <= 199;
                X_25 <= 20;
                X_26 <= 237;
                X_27 <= 198;
                X_28 <= 124;
                X_29 <= 111;
                X_30 <= 114;
                X_31 <= 78;
                X_32 <= 130;
                X_33 <= 130;
                X_34 <= 209;
                X_35 <= 203;
                X_36 <= 164;
                X_37 <= 96;
                X_38 <= 207;
                X_39 <= 136;
                X_40 <= 89;
                X_41 <= 240;
                X_42 <= 224;
                X_43 <= 140;
                X_44 <= 159;
                X_45 <= 150;
                X_46 <= 53;
                X_47 <= 77;
                X_48 <= 120;
                X_49 <= 59;
                X_50 <= 216;
                X_51 <= 49;
                X_52 <= 57;
                X_53 <= 43;
                X_54 <= 58;
                X_55 <= 111;
                out <= 0;
            end else if (number == 4) begin
                X_1 <= 122;
                X_2 <= 149;
                X_3 <= 54;
                X_4 <= 149;
                X_5 <= 199;
                X_6 <= 25;
                X_7 <= 203;
                X_8 <= 217;
                X_9 <= 175;
                X_10 <= 184;
                X_11 <= 150;
                X_12 <= 40;
                X_13 <= 163;
                X_14 <= 12;
                X_15 <= 254;
                X_16 <= 226;
                X_17 <= 170;
                X_18 <= 132;
                X_19 <= 125;
                X_20 <= 38;
                X_21 <= 234;
                X_22 <= 92;
                X_23 <= 136;
                X_24 <= 5;
                X_25 <= 153;
                X_26 <= 80;
                X_27 <= 121;
                X_28 <= 60;
                X_29 <= 189;
                X_30 <= 181;
                X_31 <= 176;
                X_32 <= 174;
                X_33 <= 78;
                X_34 <= 149;
                X_35 <= 169;
                X_36 <= 101;
                X_37 <= 113;
                X_38 <= 31;
                X_39 <= 42;
                X_40 <= 154;
                X_41 <= 136;
                X_42 <= 10;
                X_43 <= 137;
                X_44 <= 183;
                X_45 <= 115;
                X_46 <= 252;
                X_47 <= 78;
                X_48 <= 169;
                X_49 <= 236;
                X_50 <= 180;
                X_51 <= 69;
                X_52 <= 140;
                X_53 <= 153;
                X_54 <= 40;
                X_55 <= 105;
                out <= 0;  
            end else if (number == 5) begin
                X_1 <= 29;
                X_2 <= 19;
                X_3 <= 69;
                X_4 <= 74;
                X_5 <= 61;
                X_6 <= 146;
                X_7 <= 45;
                X_8 <= 255;
                X_9 <= 218;
                X_10 <= 222;
                X_11 <= 217;
                X_12 <= 135;
                X_13 <= 39;
                X_14 <= 104;
                X_15 <= 113;
                X_16 <= 39;
                X_17 <= 35;
                X_18 <= 220;
                X_19 <= 38;
                X_20 <= 14;
                X_21 <= 233;
                X_22 <= 169;
                X_23 <= 187;
                X_24 <= 166;
                X_25 <= 61;
                X_26 <= 166;
                X_27 <= 129;
                X_28 <= 121;
                X_29 <= 228;
                X_30 <= 127;
                X_31 <= 64;
                X_32 <= 22;
                X_33 <= 192;
                X_34 <= 71;
                X_35 <= 195;
                X_36 <= 189;
                X_37 <= 142;
                X_38 <= 174;
                X_39 <= 41;
                X_40 <= 189;
                X_41 <= 2;
                X_42 <= 103;
                X_43 <= 190;
                X_44 <= 166;
                X_45 <= 157;
                X_46 <= 29;
                X_47 <= 134;
                X_48 <= 242;
                X_49 <= 199;
                X_50 <= 97;
                X_51 <= 107;
                X_52 <= 51;
                X_53 <= 124;
                X_54 <= 122;
                X_55 <= 136;
                out <= 0;   
            end else if (number == 6) begin
                X_1 <= 52;
                X_2 <= 101;
                X_3 <= 61;
                X_4 <= 70;
                X_5 <= 242;
                X_6 <= 206;
                X_7 <= 223;
                X_8 <= 243;
                X_9 <= 6;
                X_10 <= 56;
                X_11 <= 192;
                X_12 <= 104;
                X_13 <= 178;
                X_14 <= 244;
                X_15 <= 4;
                X_16 <= 200;
                X_17 <= 19;
                X_18 <= 187;
                X_19 <= 238;
                X_20 <= 39;
                X_21 <= 12;
                X_22 <= 3;
                X_23 <= 102;
                X_24 <= 47;
                X_25 <= 161;
                X_26 <= 65;
                X_27 <= 163;
                X_28 <= 230;
                X_29 <= 146;
                X_30 <= 39;
                X_31 <= 139;
                X_32 <= 13;
                X_33 <= 100;
                X_34 <= 24;
                X_35 <= 38;
                X_36 <= 172;
                X_37 <= 138;
                X_38 <= 246;
                X_39 <= 93;
                X_40 <= 155;
                X_41 <= 234;
                X_42 <= 204;
                X_43 <= 213;
                X_44 <= 120;
                X_45 <= 37;
                X_46 <= 240;
                X_47 <= 174;
                X_48 <= 172;
                X_49 <= 126;
                X_50 <= 222;
                X_51 <= 24;
                X_52 <= 224;
                X_53 <= 139;
                X_54 <= 23;
                X_55 <= 241;
                out <= 0;   
            end else begin
                X_1 <= 236;
                X_2 <= 184;
                X_3 <= 170;
                X_4 <= 59;
                X_5 <= 95;
                X_6 <= 72;
                X_7 <= 210;
                X_8 <= 119;
                X_9 <= 219;
                X_10 <= 230;
                X_11 <= 74;
                X_12 <= 107;
                X_13 <= 160;
                X_14 <= 44;
                X_15 <= 131;
                X_16 <= 190;
                X_17 <= 246;
                X_18 <= 6;
                X_19 <= 121;
                X_20 <= 76;
                X_21 <= 5;
                X_22 <= 144;
                X_23 <= 193;
                X_24 <= 84;
                X_25 <= 12;
                X_26 <= 255;
                X_27 <= 107;
                X_28 <= 41;
                X_29 <= 43;
                X_30 <= 134;
                X_31 <= 228;
                X_32 <= 134;
                X_33 <= 157;
                X_34 <= 219;
                X_35 <= 106;
                X_36 <= 45;
                X_37 <= 192;
                X_38 <= 142;
                X_39 <= 218;
                X_40 <= 193;
                X_41 <= 173;
                X_42 <= 23;
                X_43 <= 163;
                X_44 <= 63;
                X_45 <= 133;
                X_46 <= 216;
                X_47 <= 60;
                X_48 <= 184;
                X_49 <= 147;
                X_50 <= 129;
                X_51 <= 133;
                X_52 <= 241;
                X_53 <= 63;
                X_54 <= 243;
                X_55 <= 22;
                out <= 0;                                                            
            end
            
        end else begin
            if (X_55 >= X_24) begin
                X_1 <= X_55 - X_24;
            end else begin
                X_1 <= X_55 - X_24 + 256;
            end
            X_55 <= X_54;
            X_54 <= X_53;
            X_53 <= X_52;
            X_52 <= X_51;
            X_51 <= X_50;
            X_50 <= X_49;
            X_49 <= X_48;
            X_48 <= X_47;
            X_47 <= X_46;
            X_46 <= X_45;
            X_45 <= X_44;
            X_44 <= X_43;
            X_43 <= X_42;
            X_42 <= X_41;
            X_41 <= X_40;
            X_40 <= X_39;
            X_39 <= X_38;
            X_38 <= X_37;
            X_37 <= X_36;
            X_36 <= X_35;
            X_35 <= X_34;
            X_34 <= X_33;
            X_33 <= X_32;
            X_32 <= X_31;
            X_31 <= X_30;
            X_30 <= X_29;
            X_29 <= X_28;
            X_28 <= X_27;
            X_27 <= X_26;
            X_26 <= X_25;
            X_25 <= X_24;
            X_24 <= X_23;
            X_23 <= X_22;
            X_22 <= X_21;
            X_21 <= X_20;
            X_20 <= X_19;
            X_19 <= X_18;
            X_18 <= X_17;
            X_17 <= X_16;
            X_16 <= X_15;
            X_15 <= X_14;
            X_14 <= X_13;
            X_13 <= X_12;
            X_12 <= X_11;
            X_11 <= X_10;
            X_10 <= X_9;
            X_9 <= X_8;
            X_8 <= X_7;
            X_7 <= X_6;
            X_6 <= X_5;
            X_5 <= X_4;
            X_4 <= X_3;
            X_3 <= X_2;
            X_2 <= X_1;
            out <= X_1;      
        end
    end
endmodule
