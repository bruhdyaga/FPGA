`timescale 1ns/10ps

module channel_cmplx_table (
		clk,
		reset_n,
		adc_re,
		adc_im,
		cos_product,
		sin_product,		
		phase_addr,
		cmplx_product_re,
		cmplx_product_im
		);
    
	input clk;
	input reset_n;
	input [1 : 0] adc_re;
	input [1 : 0] adc_im;
	input signed [4 : 0] cos_product;
	input signed [4 : 0] sin_product;
	input [4 : 0] phase_addr;
	output signed [4 : 0] cmplx_product_re;
	output signed [4 : 0] cmplx_product_im;
	    
	reg  signed [4 : 0] cos_product_r;
	reg  signed [4 : 0] sin_product_r;
	reg  signed [5 : 0] cmplx_product_r;
	reg  signed [4 : 0] cmplx_product_c;
	wire signed [5:0] cmplx_product_re_wide;
	wire signed [6:0] cmplx_product_im_wide;
    
	always @(*) begin
		case ({adc_re[1 : 0], adc_im[1 : 0], phase_addr[4 : 0]})
			{2'b00, 2'b00, 5'd0}     : cmplx_product_c = 5'h3;
			{2'b00, 2'b00, 5'd1}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b00, 5'd2}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b00, 5'd3}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b00, 5'd4}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b00, 5'd5}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b00, 5'd6}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b00, 5'd7}     : cmplx_product_c = 5'h3;
			{2'b00, 2'b00, 5'd8}     : cmplx_product_c = 5'h3;
			{2'b00, 2'b00, 5'd9}     : cmplx_product_c = 5'h2;
			{2'b00, 2'b00, 5'd10}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b00, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b00, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b00, 5'd13}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b00, 5'd14}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b00, 5'd15}    : cmplx_product_c = 5'h1d;			
			{2'b00, 2'b00, 5'd16}    : cmplx_product_c = 5'h1d;
			{2'b00, 2'b00, 5'd17}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b00, 5'd18}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b00, 5'd19}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b00, 5'd20}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b00, 5'd21}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b00, 5'd22}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b00, 5'd23}    : cmplx_product_c = 5'h1d;
			{2'b00, 2'b00, 5'd24}    : cmplx_product_c = 5'h1d;
			{2'b00, 2'b00, 5'd25}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b00, 5'd26}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b00, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b00, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b00, 5'd29}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b00, 5'd30}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b00, 5'd31}    : cmplx_product_c = 5'h3;
			
			{2'b00, 2'b01, 5'd0}     : cmplx_product_c = 5'h6;
			{2'b00, 2'b01, 5'd1}     : cmplx_product_c = 5'h8;
			{2'b00, 2'b01, 5'd2}     : cmplx_product_c = 5'h8;
			{2'b00, 2'b01, 5'd3}     : cmplx_product_c = 5'h8;
			{2'b00, 2'b01, 5'd4}     : cmplx_product_c = 5'h8;
			{2'b00, 2'b01, 5'd5}     : cmplx_product_c = 5'h8;
			{2'b00, 2'b01, 5'd6}     : cmplx_product_c = 5'h8;
			{2'b00, 2'b01, 5'd7}     : cmplx_product_c = 5'h6;
			{2'b00, 2'b01, 5'd8}     : cmplx_product_c = 5'h6;
			{2'b00, 2'b01, 5'd9}     : cmplx_product_c = 5'h4;
			{2'b00, 2'b01, 5'd10}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b01, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b01, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b01, 5'd13}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b01, 5'd14}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b01, 5'd15}    : cmplx_product_c = 5'h1a;			
			{2'b00, 2'b01, 5'd16}    : cmplx_product_c = 5'h1a;
			{2'b00, 2'b01, 5'd17}    : cmplx_product_c = 5'h18;
			{2'b00, 2'b01, 5'd18}    : cmplx_product_c = 5'h18;
			{2'b00, 2'b01, 5'd19}    : cmplx_product_c = 5'h18;
			{2'b00, 2'b01, 5'd20}    : cmplx_product_c = 5'h18;
			{2'b00, 2'b01, 5'd21}    : cmplx_product_c = 5'h18;
			{2'b00, 2'b01, 5'd22}    : cmplx_product_c = 5'h18;
			{2'b00, 2'b01, 5'd23}    : cmplx_product_c = 5'h1a;
			{2'b00, 2'b01, 5'd24}    : cmplx_product_c = 5'h1a;
			{2'b00, 2'b01, 5'd25}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b01, 5'd26}    : cmplx_product_c = 5'h1c;
			{2'b00, 2'b01, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b01, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b01, 5'd29}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b01, 5'd30}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b01, 5'd31}    : cmplx_product_c = 5'h6;
			
			{2'b00, 2'b10, 5'd0}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd1}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd2}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd3}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd4}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd5}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd6}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd7}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd8}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd9}     : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd10}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd13}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd14}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd15}    : cmplx_product_c = 5'h0;			
			{2'b00, 2'b10, 5'd16}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd17}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd18}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd19}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd20}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd21}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd22}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd23}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd24}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd25}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd26}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd29}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd30}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b10, 5'd31}    : cmplx_product_c = 5'h0;
			
			{2'b00, 2'b11, 5'd0}     : cmplx_product_c = 5'h1d;
			{2'b00, 2'b11, 5'd1}     : cmplx_product_c = 5'h1c;
			{2'b00, 2'b11, 5'd2}     : cmplx_product_c = 5'h1c;
			{2'b00, 2'b11, 5'd3}     : cmplx_product_c = 5'h1c;
			{2'b00, 2'b11, 5'd4}     : cmplx_product_c = 5'h1c;
			{2'b00, 2'b11, 5'd5}     : cmplx_product_c = 5'h1c;
			{2'b00, 2'b11, 5'd6}     : cmplx_product_c = 5'h1c;
			{2'b00, 2'b11, 5'd7}     : cmplx_product_c = 5'h1d;
			{2'b00, 2'b11, 5'd8}     : cmplx_product_c = 5'h1d;
			{2'b00, 2'b11, 5'd9}     : cmplx_product_c = 5'h1e;
			{2'b00, 2'b11, 5'd10}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b11, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b11, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b11, 5'd13}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b11, 5'd14}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b11, 5'd15}    : cmplx_product_c = 5'h3;			
			{2'b00, 2'b11, 5'd16}    : cmplx_product_c = 5'h3;
			{2'b00, 2'b11, 5'd17}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b11, 5'd18}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b11, 5'd19}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b11, 5'd20}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b11, 5'd21}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b11, 5'd22}    : cmplx_product_c = 5'h4;
			{2'b00, 2'b11, 5'd23}    : cmplx_product_c = 5'h3;
			{2'b00, 2'b11, 5'd24}    : cmplx_product_c = 5'h3;
			{2'b00, 2'b11, 5'd25}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b11, 5'd26}    : cmplx_product_c = 5'h2;
			{2'b00, 2'b11, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b11, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b00, 2'b11, 5'd29}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b11, 5'd30}    : cmplx_product_c = 5'h1e;
			{2'b00, 2'b11, 5'd31}    : cmplx_product_c = 5'h1d;
			
			{2'b01, 2'b00, 5'd0}     : cmplx_product_c = 5'h6;
			{2'b01, 2'b00, 5'd1}     : cmplx_product_c = 5'h8;
			{2'b01, 2'b00, 5'd2}     : cmplx_product_c = 5'h8;
			{2'b01, 2'b00, 5'd3}     : cmplx_product_c = 5'h8;
			{2'b01, 2'b00, 5'd4}     : cmplx_product_c = 5'h8;
			{2'b01, 2'b00, 5'd5}     : cmplx_product_c = 5'h8;
			{2'b01, 2'b00, 5'd6}     : cmplx_product_c = 5'h8;
			{2'b01, 2'b00, 5'd7}     : cmplx_product_c = 5'h6;
			{2'b01, 2'b00, 5'd8}     : cmplx_product_c = 5'h6;
			{2'b01, 2'b00, 5'd9}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b00, 5'd10}    : cmplx_product_c = 5'h4;
			{2'b01, 2'b00, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b00, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b00, 5'd13}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b00, 5'd14}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b00, 5'd15}    : cmplx_product_c = 5'h1a;			
			{2'b01, 2'b00, 5'd16}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b00, 5'd17}    : cmplx_product_c = 5'h18;
			{2'b01, 2'b00, 5'd18}    : cmplx_product_c = 5'h18;
			{2'b01, 2'b00, 5'd19}    : cmplx_product_c = 5'h18;
			{2'b01, 2'b00, 5'd20}    : cmplx_product_c = 5'h18;
			{2'b01, 2'b00, 5'd21}    : cmplx_product_c = 5'h18;
			{2'b01, 2'b00, 5'd22}    : cmplx_product_c = 5'h18;
			{2'b01, 2'b00, 5'd23}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b00, 5'd24}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b00, 5'd25}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b00, 5'd26}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b00, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b00, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b00, 5'd29}    : cmplx_product_c = 5'h4;
			{2'b01, 2'b00, 5'd30}    : cmplx_product_c = 5'h4;
			{2'b01, 2'b00, 5'd31}    : cmplx_product_c = 5'h6;
			
			{2'b01, 2'b01, 5'd0}     : cmplx_product_c = 5'h9;
			{2'b01, 2'b01, 5'd1}     : cmplx_product_c = 5'hc;
			{2'b01, 2'b01, 5'd2}     : cmplx_product_c = 5'hc;
			{2'b01, 2'b01, 5'd3}     : cmplx_product_c = 5'hc;
			{2'b01, 2'b01, 5'd4}     : cmplx_product_c = 5'hc;
			{2'b01, 2'b01, 5'd5}     : cmplx_product_c = 5'hc;
			{2'b01, 2'b01, 5'd6}     : cmplx_product_c = 5'hc;
			{2'b01, 2'b01, 5'd7}     : cmplx_product_c = 5'h9;
			{2'b01, 2'b01, 5'd8}     : cmplx_product_c = 5'h9;
			{2'b01, 2'b01, 5'd9}     : cmplx_product_c = 5'h6;
			{2'b01, 2'b01, 5'd10}    : cmplx_product_c = 5'h6;
			{2'b01, 2'b01, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b01, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b01, 5'd13}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b01, 5'd14}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b01, 5'd15}    : cmplx_product_c = 5'h17;			
			{2'b01, 2'b01, 5'd16}    : cmplx_product_c = 5'h17;
			{2'b01, 2'b01, 5'd17}    : cmplx_product_c = 5'h14;
			{2'b01, 2'b01, 5'd18}    : cmplx_product_c = 5'h14;
			{2'b01, 2'b01, 5'd19}    : cmplx_product_c = 5'h14;
			{2'b01, 2'b01, 5'd20}    : cmplx_product_c = 5'h14;
			{2'b01, 2'b01, 5'd21}    : cmplx_product_c = 5'h14;
			{2'b01, 2'b01, 5'd22}    : cmplx_product_c = 5'h14;
			{2'b01, 2'b01, 5'd23}    : cmplx_product_c = 5'h17;
			{2'b01, 2'b01, 5'd24}    : cmplx_product_c = 5'h17;
			{2'b01, 2'b01, 5'd25}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b01, 5'd26}    : cmplx_product_c = 5'h1a;
			{2'b01, 2'b01, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b01, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b01, 5'd29}    : cmplx_product_c = 5'h6;
			{2'b01, 2'b01, 5'd30}    : cmplx_product_c = 5'h6;
			{2'b01, 2'b01, 5'd31}    : cmplx_product_c = 5'h9;
			
			{2'b01, 2'b10, 5'd0}     : cmplx_product_c = 5'h3;
			{2'b01, 2'b10, 5'd1}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b10, 5'd2}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b10, 5'd3}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b10, 5'd4}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b10, 5'd5}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b10, 5'd6}     : cmplx_product_c = 5'h4;
			{2'b01, 2'b10, 5'd7}     : cmplx_product_c = 5'h3;
			{2'b01, 2'b10, 5'd8}     : cmplx_product_c = 5'h3;
			{2'b01, 2'b10, 5'd9}     : cmplx_product_c = 5'h2;
			{2'b01, 2'b10, 5'd10}    : cmplx_product_c = 5'h2;
			{2'b01, 2'b10, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b10, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b10, 5'd13}    : cmplx_product_c = 5'h1e;
			{2'b01, 2'b10, 5'd14}    : cmplx_product_c = 5'h1e;
			{2'b01, 2'b10, 5'd15}    : cmplx_product_c = 5'h1d;			
			{2'b01, 2'b10, 5'd16}    : cmplx_product_c = 5'h1d;
			{2'b01, 2'b10, 5'd17}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b10, 5'd18}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b10, 5'd19}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b10, 5'd20}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b10, 5'd21}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b10, 5'd22}    : cmplx_product_c = 5'h1c;
			{2'b01, 2'b10, 5'd23}    : cmplx_product_c = 5'h1d;
			{2'b01, 2'b10, 5'd24}    : cmplx_product_c = 5'h1d;
			{2'b01, 2'b10, 5'd25}    : cmplx_product_c = 5'h1e;
			{2'b01, 2'b10, 5'd26}    : cmplx_product_c = 5'h1e;
			{2'b01, 2'b10, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b10, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b10, 5'd29}    : cmplx_product_c = 5'h2;
			{2'b01, 2'b10, 5'd30}    : cmplx_product_c = 5'h2;
			{2'b01, 2'b10, 5'd31}    : cmplx_product_c = 5'h3;
			
			{2'b01, 2'b11, 5'd0}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd1}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd2}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd3}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd4}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd5}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd6}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd7}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd8}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd9}     : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd10}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd13}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd14}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd15}    : cmplx_product_c = 5'h0;			
			{2'b01, 2'b11, 5'd16}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd17}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd18}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd19}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd20}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd21}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd22}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd23}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd24}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd25}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd26}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd29}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd30}    : cmplx_product_c = 5'h0;
			{2'b01, 2'b11, 5'd31}    : cmplx_product_c = 5'h0;
			
			{2'b10, 2'b00, 5'd0}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd1}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd2}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd3}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd4}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd5}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd6}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd7}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd8}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd9}     : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd10}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd13}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd14}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd15}    : cmplx_product_c = 5'h0;			
			{2'b10, 2'b00, 5'd16}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd17}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd18}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd19}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd20}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd21}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd22}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd23}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd24}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd25}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd26}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd29}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd30}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b00, 5'd31}    : cmplx_product_c = 5'h0;
			
			{2'b10, 2'b01, 5'd0}     : cmplx_product_c = 5'h1d;
			{2'b10, 2'b01, 5'd1}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b01, 5'd2}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b01, 5'd3}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b01, 5'd4}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b01, 5'd5}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b01, 5'd6}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b01, 5'd7}     : cmplx_product_c = 5'h1d;
			{2'b10, 2'b01, 5'd8}     : cmplx_product_c = 5'h1d;
			{2'b10, 2'b01, 5'd9}     : cmplx_product_c = 5'h1e;
			{2'b10, 2'b01, 5'd10}    : cmplx_product_c = 5'h1e;
			{2'b10, 2'b01, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b01, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b01, 5'd13}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b01, 5'd14}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b01, 5'd15}    : cmplx_product_c = 5'h3;			
			{2'b10, 2'b01, 5'd16}    : cmplx_product_c = 5'h3;
			{2'b10, 2'b01, 5'd17}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b01, 5'd18}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b01, 5'd19}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b01, 5'd20}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b01, 5'd21}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b01, 5'd22}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b01, 5'd23}    : cmplx_product_c = 5'h3;
			{2'b10, 2'b01, 5'd24}    : cmplx_product_c = 5'h3;
			{2'b10, 2'b01, 5'd25}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b01, 5'd26}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b01, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b01, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b01, 5'd29}    : cmplx_product_c = 5'h1e;
			{2'b10, 2'b01, 5'd30}    : cmplx_product_c = 5'h1e;
			{2'b10, 2'b01, 5'd31}    : cmplx_product_c = 5'h1d;
			
			{2'b10, 2'b10, 5'd0}     : cmplx_product_c = 5'h1d;
			{2'b10, 2'b10, 5'd1}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b10, 5'd2}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b10, 5'd3}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b10, 5'd4}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b10, 5'd5}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b10, 5'd6}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b10, 5'd7}     : cmplx_product_c = 5'h1d;
			{2'b10, 2'b10, 5'd8}     : cmplx_product_c = 5'h1d;
			{2'b10, 2'b10, 5'd9}     : cmplx_product_c = 5'h1e;
			{2'b10, 2'b10, 5'd10}    : cmplx_product_c = 5'h1e;
			{2'b10, 2'b10, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b10, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b10, 5'd13}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b10, 5'd14}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b10, 5'd15}    : cmplx_product_c = 5'h3;			
			{2'b10, 2'b10, 5'd16}    : cmplx_product_c = 5'h3;
			{2'b10, 2'b10, 5'd17}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b10, 5'd18}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b10, 5'd19}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b10, 5'd20}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b10, 5'd21}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b10, 5'd22}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b10, 5'd23}    : cmplx_product_c = 5'h3;
			{2'b10, 2'b10, 5'd24}    : cmplx_product_c = 5'h3;
			{2'b10, 2'b10, 5'd25}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b10, 5'd26}    : cmplx_product_c = 5'h2;
			{2'b10, 2'b10, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b10, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b10, 5'd29}    : cmplx_product_c = 5'h1e;
			{2'b10, 2'b10, 5'd30}    : cmplx_product_c = 5'h1e;
			{2'b10, 2'b10, 5'd31}    : cmplx_product_c = 5'h1d;
			
			{2'b10, 2'b11, 5'd0}     : cmplx_product_c = 5'h1a;
			{2'b10, 2'b11, 5'd1}     : cmplx_product_c = 5'h18;
			{2'b10, 2'b11, 5'd2}     : cmplx_product_c = 5'h18;
			{2'b10, 2'b11, 5'd3}     : cmplx_product_c = 5'h18;
			{2'b10, 2'b11, 5'd4}     : cmplx_product_c = 5'h18;
			{2'b10, 2'b11, 5'd5}     : cmplx_product_c = 5'h18;
			{2'b10, 2'b11, 5'd6}     : cmplx_product_c = 5'h18;
			{2'b10, 2'b11, 5'd7}     : cmplx_product_c = 5'h1a;
			{2'b10, 2'b11, 5'd8}     : cmplx_product_c = 5'h1a;
			{2'b10, 2'b11, 5'd9}     : cmplx_product_c = 5'h1c;
			{2'b10, 2'b11, 5'd10}    : cmplx_product_c = 5'h1c;
			{2'b10, 2'b11, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b11, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b11, 5'd13}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b11, 5'd14}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b11, 5'd15}    : cmplx_product_c = 5'h6;			
			{2'b10, 2'b11, 5'd16}    : cmplx_product_c = 5'h6;
			{2'b10, 2'b11, 5'd17}    : cmplx_product_c = 5'h8;
			{2'b10, 2'b11, 5'd18}    : cmplx_product_c = 5'h8;
			{2'b10, 2'b11, 5'd19}    : cmplx_product_c = 5'h8;
			{2'b10, 2'b11, 5'd20}    : cmplx_product_c = 5'h8;
			{2'b10, 2'b11, 5'd21}    : cmplx_product_c = 5'h8;
			{2'b10, 2'b11, 5'd22}    : cmplx_product_c = 5'h8;
			{2'b10, 2'b11, 5'd23}    : cmplx_product_c = 5'h6;
			{2'b10, 2'b11, 5'd24}    : cmplx_product_c = 5'h6;
			{2'b10, 2'b11, 5'd25}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b11, 5'd26}    : cmplx_product_c = 5'h4;
			{2'b10, 2'b11, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b11, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b10, 2'b11, 5'd29}    : cmplx_product_c = 5'h1c;
			{2'b10, 2'b11, 5'd30}    : cmplx_product_c = 5'h1c;
			{2'b10, 2'b11, 5'd31}    : cmplx_product_c = 5'h1a;
			
			{2'b11, 2'b00, 5'd0}     : cmplx_product_c = 5'h1d;
			{2'b11, 2'b00, 5'd1}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b00, 5'd2}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b00, 5'd3}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b00, 5'd4}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b00, 5'd5}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b00, 5'd6}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b00, 5'd7}     : cmplx_product_c = 5'h1d;
			{2'b11, 2'b00, 5'd8}     : cmplx_product_c = 5'h1d;
			{2'b11, 2'b00, 5'd9}     : cmplx_product_c = 5'h1e;
			{2'b11, 2'b00, 5'd10}    : cmplx_product_c = 5'h1e;
			{2'b11, 2'b00, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b00, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b00, 5'd13}    : cmplx_product_c = 5'h2;
			{2'b11, 2'b00, 5'd14}    : cmplx_product_c = 5'h2;
			{2'b11, 2'b00, 5'd15}    : cmplx_product_c = 5'h3;			
			{2'b11, 2'b00, 5'd16}    : cmplx_product_c = 5'h3;
			{2'b11, 2'b00, 5'd17}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b00, 5'd18}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b00, 5'd19}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b00, 5'd20}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b00, 5'd21}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b00, 5'd22}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b00, 5'd23}    : cmplx_product_c = 5'h3;
			{2'b11, 2'b00, 5'd24}    : cmplx_product_c = 5'h3;
			{2'b11, 2'b00, 5'd25}    : cmplx_product_c = 5'h2;
			{2'b11, 2'b00, 5'd26}    : cmplx_product_c = 5'h2;
			{2'b11, 2'b00, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b00, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b00, 5'd29}    : cmplx_product_c = 5'h1e;
			{2'b11, 2'b00, 5'd30}    : cmplx_product_c = 5'h1e;
			{2'b11, 2'b00, 5'd31}    : cmplx_product_c = 5'h1d;
			
			{2'b11, 2'b01, 5'd0}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd1}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd2}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd3}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd4}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd5}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd6}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd7}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd8}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd9}     : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd10}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd13}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd14}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd15}    : cmplx_product_c = 5'h0;			
			{2'b11, 2'b01, 5'd16}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd17}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd18}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd19}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd20}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd21}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd22}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd23}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd24}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd25}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd26}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd29}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd30}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b01, 5'd31}    : cmplx_product_c = 5'h0;
			
			{2'b11, 2'b10, 5'd0}     : cmplx_product_c = 5'h1a;
			{2'b11, 2'b10, 5'd1}     : cmplx_product_c = 5'h18;
			{2'b11, 2'b10, 5'd2}     : cmplx_product_c = 5'h18;
			{2'b11, 2'b10, 5'd3}     : cmplx_product_c = 5'h18;
			{2'b11, 2'b10, 5'd4}     : cmplx_product_c = 5'h18;
			{2'b11, 2'b10, 5'd5}     : cmplx_product_c = 5'h18;
			{2'b11, 2'b10, 5'd6}     : cmplx_product_c = 5'h18;
			{2'b11, 2'b10, 5'd7}     : cmplx_product_c = 5'h1a;
			{2'b11, 2'b10, 5'd8}     : cmplx_product_c = 5'h1a;
			{2'b11, 2'b10, 5'd9}     : cmplx_product_c = 5'h1c;
			{2'b11, 2'b10, 5'd10}    : cmplx_product_c = 5'h1c;
			{2'b11, 2'b10, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b10, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b10, 5'd13}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b10, 5'd14}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b10, 5'd15}    : cmplx_product_c = 5'h6;			
			{2'b11, 2'b10, 5'd16}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b10, 5'd17}    : cmplx_product_c = 5'h8;
			{2'b11, 2'b10, 5'd18}    : cmplx_product_c = 5'h8;
			{2'b11, 2'b10, 5'd19}    : cmplx_product_c = 5'h8;
			{2'b11, 2'b10, 5'd20}    : cmplx_product_c = 5'h8;
			{2'b11, 2'b10, 5'd21}    : cmplx_product_c = 5'h8;
			{2'b11, 2'b10, 5'd22}    : cmplx_product_c = 5'h8;
			{2'b11, 2'b10, 5'd23}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b10, 5'd24}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b10, 5'd25}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b10, 5'd26}    : cmplx_product_c = 5'h4;
			{2'b11, 2'b10, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b10, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b10, 5'd29}    : cmplx_product_c = 5'h1c;
			{2'b11, 2'b10, 5'd30}    : cmplx_product_c = 5'h1c;
			{2'b11, 2'b10, 5'd31}    : cmplx_product_c = 5'h1a;
			
			{2'b11, 2'b11, 5'd0}     : cmplx_product_c = 5'h17;
			{2'b11, 2'b11, 5'd1}     : cmplx_product_c = 5'h14;
			{2'b11, 2'b11, 5'd2}     : cmplx_product_c = 5'h14;
			{2'b11, 2'b11, 5'd3}     : cmplx_product_c = 5'h14;
			{2'b11, 2'b11, 5'd4}     : cmplx_product_c = 5'h14;
			{2'b11, 2'b11, 5'd5}     : cmplx_product_c = 5'h14;
			{2'b11, 2'b11, 5'd6}     : cmplx_product_c = 5'h14;
			{2'b11, 2'b11, 5'd7}     : cmplx_product_c = 5'h17;
			{2'b11, 2'b11, 5'd8}     : cmplx_product_c = 5'h17;
			{2'b11, 2'b11, 5'd9}     : cmplx_product_c = 5'h1a;
			{2'b11, 2'b11, 5'd10}    : cmplx_product_c = 5'h1a;
			{2'b11, 2'b11, 5'd11}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b11, 5'd12}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b11, 5'd13}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b11, 5'd14}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b11, 5'd15}    : cmplx_product_c = 5'h9;			
			{2'b11, 2'b11, 5'd16}    : cmplx_product_c = 5'h9;
			{2'b11, 2'b11, 5'd17}    : cmplx_product_c = 5'hc;
			{2'b11, 2'b11, 5'd18}    : cmplx_product_c = 5'hc;
			{2'b11, 2'b11, 5'd19}    : cmplx_product_c = 5'hc;
			{2'b11, 2'b11, 5'd20}    : cmplx_product_c = 5'hc;
			{2'b11, 2'b11, 5'd21}    : cmplx_product_c = 5'hc;
			{2'b11, 2'b11, 5'd22}    : cmplx_product_c = 5'hc;
			{2'b11, 2'b11, 5'd23}    : cmplx_product_c = 5'h9;
			{2'b11, 2'b11, 5'd24}    : cmplx_product_c = 5'h9;
			{2'b11, 2'b11, 5'd25}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b11, 5'd26}    : cmplx_product_c = 5'h6;
			{2'b11, 2'b11, 5'd27}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b11, 5'd28}    : cmplx_product_c = 5'h0;
			{2'b11, 2'b11, 5'd29}    : cmplx_product_c = 5'h1a;
			{2'b11, 2'b11, 5'd30}    : cmplx_product_c = 5'h1a;
			{2'b11, 2'b11, 5'd31}    : cmplx_product_c = 5'h17;		
		endcase
	end
	
	always @ (posedge clk or negedge reset_n) begin
        if (reset_n == 1'b0) begin
            cos_product_r <= 5'b0;
        	sin_product_r <= 5'b0;
            cmplx_product_r <= 6'b0;
        end
        else begin
        	cos_product_r <= cos_product;
            sin_product_r <= sin_product;
            cmplx_product_r <= cmplx_product_c <<< 1;
        end
    end
    assign cmplx_product_re_wide = $signed(cos_product_r - sin_product_r);
    assign cmplx_product_re = cmplx_product_re_wide[5:1];
	assign cmplx_product_im_wide = $signed(cmplx_product_r - cos_product_r - sin_product_r);
    assign cmplx_product_im = cmplx_product_im_wide[5:1];
    

endmodule
