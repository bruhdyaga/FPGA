module randn_u#(
    parameter number = 0 // Порядковый номер блока (отличаются зерном)
)
(
    input                     clk,
    input                     set,
    output logic signed [7:0] out
);

logic signed [7:0] X [55:1];

generate
always_ff@(posedge clk)
if(set) begin
    if(number == 0) begin
        X[1]  <= 208;
        X[2]  <= 231;
        X[3]  <= 32;
        X[4]  <= 233;
        X[5]  <= 161;
        X[6]  <= 24;
        X[7]  <= 71;
        X[8]  <= 140;
        X[9]  <= 245;
        X[10] <= 247;
        X[11] <= 40;
        X[12] <= 248;
        X[13] <= 245;
        X[14] <= 124;
        X[15] <= 204;
        X[16] <= 36;
        X[17] <= 107;
        X[18] <= 234;
        X[19] <= 202;
        X[20] <= 245;
        X[21] <= 167;
        X[22] <= 9;
        X[23] <= 217;
        X[24] <= 239;
        X[25] <= 173;
        X[26] <= 193;
        X[27] <= 190;
        X[28] <= 100;
        X[29] <= 167;
        X[30] <= 43;
        X[31] <= 180;
        X[32] <= 8;
        X[33] <= 70;
        X[34] <= 11;
        X[35] <= 24;
        X[36] <= 210;
        X[37] <= 177;
        X[38] <= 81;
        X[39] <= 243;
        X[40] <= 8;
        X[41] <= 112;
        X[42] <= 97;
        X[43] <= 195;
        X[44] <= 203;
        X[45] <= 47;
        X[46] <= 125;
        X[47] <= 114;
        X[48] <= 165;
        X[49] <= 181;
        X[50] <= 193;
        X[51] <= 70;
        X[52] <= 174;
        X[53] <= 167;
        X[54] <= 41;
        X[55] <= 30;
        out   <= 0;
    end else if (number == 1) begin
        X[1]  <= 127;
        X[2]  <= 245;
        X[3]  <= 87;
        X[4]  <= 149;
        X[5]  <= 57;
        X[6]  <= 192;
        X[7]  <= 65;
        X[8]  <= 129;
        X[9]  <= 178;
        X[10] <= 228;
        X[11] <= 245;
        X[12] <= 140;
        X[13] <= 35;
        X[14] <= 38;
        X[15] <= 65;
        X[16] <= 215;
        X[17] <= 65;
        X[18] <= 208;
        X[19] <= 62;
        X[20] <= 237;
        X[21] <= 89;
        X[22] <= 50;
        X[23] <= 64;
        X[24] <= 157;
        X[25] <= 121;
        X[26] <= 90;
        X[27] <= 212;
        X[28] <= 149;
        X[29] <= 140;
        X[30] <= 234;
        X[31] <= 73;
        X[32] <= 193;
        X[33] <= 192;
        X[34] <= 97;
        X[35] <= 145;
        X[36] <= 19;
        X[37] <= 13;
        X[38] <= 135;
        X[39] <= 199;
        X[40] <= 239;
        X[41] <= 33;
        X[42] <= 145;
        X[43] <= 120;
        X[44] <= 3;
        X[45] <= 86;
        X[46] <= 41;
        X[47] <= 203;
        X[48] <= 79;
        X[49] <= 135;
        X[50] <= 42;
        X[51] <= 154;
        X[52] <= 67;
        X[53] <= 167;
        X[54] <= 176;
        X[55] <= 191;
        out   <= 0;
    end else if (number == 2) begin
        X[1]  <= 115;
        X[2]  <= 21;
        X[3]  <= 58;
        X[4]  <= 233;
        X[5]  <= 39;
        X[6]  <= 211;
        X[7]  <= 137;
        X[8]  <= 255;
        X[9]  <= 20;
        X[10] <= 113;
        X[11] <= 27;
        X[12] <= 246;
        X[13] <= 1;
        X[14] <= 198;
        X[15] <= 209;
        X[16] <= 222;
        X[17] <= 21;
        X[18] <= 102;
        X[19] <= 66;
        X[20] <= 204;
        X[21] <= 110;
        X[22] <= 233;
        X[23] <= 46;
        X[24] <= 67;
        X[25] <= 37;
        X[26] <= 34;
        X[27] <= 222;
        X[28] <= 148;
        X[29] <= 140;
        X[30] <= 37;
        X[31] <= 218;
        X[32] <= 159;
        X[33] <= 89;
        X[34] <= 131;
        X[35] <= 102;
        X[36] <= 19;
        X[37] <= 61;
        X[38] <= 31;
        X[39] <= 47;
        X[40] <= 61;
        X[41] <= 106;
        X[42] <= 12;
        X[43] <= 231;
        X[44] <= 241;
        X[45] <= 125;
        X[46] <= 125;
        X[47] <= 86;
        X[48] <= 230;
        X[49] <= 94;
        X[50] <= 28;
        X[51] <= 199;
        X[52] <= 99;
        X[53] <= 61;
        X[54] <= 103;
        X[55] <= 24;
        out   <= 0;
    end else if (number == 3) begin
        X[1]  <= 33;
        X[2]  <= 241;
        X[3]  <= 244;
        X[4]  <= 147;
        X[5]  <= 15;
        X[6]  <= 60;
        X[7]  <= 90;
        X[8]  <= 210;
        X[9]  <= 3;
        X[10] <= 11;
        X[11] <= 43;
        X[12] <= 166;
        X[13] <= 187;
        X[14] <= 165;
        X[15] <= 115;
        X[16] <= 140;
        X[17] <= 75;
        X[18] <= 190;
        X[19] <= 48;
        X[20] <= 175;
        X[21] <= 46;
        X[22] <= 94;
        X[23] <= 160;
        X[24] <= 199;
        X[25] <= 20;
        X[26] <= 237;
        X[27] <= 198;
        X[28] <= 124;
        X[29] <= 111;
        X[30] <= 114;
        X[31] <= 78;
        X[32] <= 130;
        X[33] <= 130;
        X[34] <= 209;
        X[35] <= 203;
        X[36] <= 164;
        X[37] <= 96;
        X[38] <= 207;
        X[39] <= 136;
        X[40] <= 89;
        X[41] <= 240;
        X[42] <= 224;
        X[43] <= 140;
        X[44] <= 159;
        X[45] <= 150;
        X[46] <= 53;
        X[47] <= 77;
        X[48] <= 120;
        X[49] <= 59;
        X[50] <= 216;
        X[51] <= 49;
        X[52] <= 57;
        X[53] <= 43;
        X[54] <= 58;
        X[55] <= 111;
        out   <= 0;
    end else if (number == 4) begin
        X[1]  <= 122;
        X[2]  <= 149;
        X[3]  <= 54;
        X[4]  <= 149;
        X[5]  <= 199;
        X[6]  <= 25;
        X[7]  <= 203;
        X[8]  <= 217;
        X[9]  <= 175;
        X[10] <= 184;
        X[11] <= 150;
        X[12] <= 40;
        X[13] <= 163;
        X[14] <= 12;
        X[15] <= 254;
        X[16] <= 226;
        X[17] <= 170;
        X[18] <= 132;
        X[19] <= 125;
        X[20] <= 38;
        X[21] <= 234;
        X[22] <= 92;
        X[23] <= 136;
        X[24] <= 5;
        X[25] <= 153;
        X[26] <= 80;
        X[27] <= 121;
        X[28] <= 60;
        X[29] <= 189;
        X[30] <= 181;
        X[31] <= 176;
        X[32] <= 174;
        X[33] <= 78;
        X[34] <= 149;
        X[35] <= 169;
        X[36] <= 101;
        X[37] <= 113;
        X[38] <= 31;
        X[39] <= 42;
        X[40] <= 154;
        X[41] <= 136;
        X[42] <= 10;
        X[43] <= 137;
        X[44] <= 183;
        X[45] <= 115;
        X[46] <= 252;
        X[47] <= 78;
        X[48] <= 169;
        X[49] <= 236;
        X[50] <= 180;
        X[51] <= 69;
        X[52] <= 140;
        X[53] <= 153;
        X[54] <= 40;
        X[55] <= 105;
        out   <= 0;
    end else if (number == 5) begin
        X[1]  <= 29;
        X[2]  <= 19;
        X[3]  <= 69;
        X[4]  <= 74;
        X[5]  <= 61;
        X[6]  <= 146;
        X[7]  <= 45;
        X[8]  <= 255;
        X[9]  <= 218;
        X[10] <= 222;
        X[11] <= 217;
        X[12] <= 135;
        X[13] <= 39;
        X[14] <= 104;
        X[15] <= 113;
        X[16] <= 39;
        X[17] <= 35;
        X[18] <= 220;
        X[19] <= 38;
        X[20] <= 14;
        X[21] <= 233;
        X[22] <= 169;
        X[23] <= 187;
        X[24] <= 166;
        X[25] <= 61;
        X[26] <= 166;
        X[27] <= 129;
        X[28] <= 121;
        X[29] <= 228;
        X[30] <= 127;
        X[31] <= 64;
        X[32] <= 22;
        X[33] <= 192;
        X[34] <= 71;
        X[35] <= 195;
        X[36] <= 189;
        X[37] <= 142;
        X[38] <= 174;
        X[39] <= 41;
        X[40] <= 189;
        X[41] <= 2;
        X[42] <= 103;
        X[43] <= 190;
        X[44] <= 166;
        X[45] <= 157;
        X[46] <= 29;
        X[47] <= 134;
        X[48] <= 242;
        X[49] <= 199;
        X[50] <= 97;
        X[51] <= 107;
        X[52] <= 51;
        X[53] <= 124;
        X[54] <= 122;
        X[55] <= 136;
        out   <= 0;
    end else if (number == 6) begin
        X[1]  <= 52;
        X[2]  <= 101;
        X[3]  <= 61;
        X[4]  <= 70;
        X[5]  <= 242;
        X[6]  <= 206;
        X[7]  <= 223;
        X[8]  <= 243;
        X[9]  <= 6;
        X[10] <= 56;
        X[11] <= 192;
        X[12] <= 104;
        X[13] <= 178;
        X[14] <= 244;
        X[15] <= 4;
        X[16] <= 200;
        X[17] <= 19;
        X[18] <= 187;
        X[19] <= 238;
        X[20] <= 39;
        X[21] <= 12;
        X[22] <= 3;
        X[23] <= 102;
        X[24] <= 47;
        X[25] <= 161;
        X[26] <= 65;
        X[27] <= 163;
        X[28] <= 230;
        X[29] <= 146;
        X[30] <= 39;
        X[31] <= 139;
        X[32] <= 13;
        X[33] <= 100;
        X[34] <= 24;
        X[35] <= 38;
        X[36] <= 172;
        X[37] <= 138;
        X[38] <= 246;
        X[39] <= 93;
        X[40] <= 155;
        X[41] <= 234;
        X[42] <= 204;
        X[43] <= 213;
        X[44] <= 120;
        X[45] <= 37;
        X[46] <= 240;
        X[47] <= 174;
        X[48] <= 172;
        X[49] <= 126;
        X[50] <= 222;
        X[51] <= 24;
        X[52] <= 224;
        X[53] <= 139;
        X[54] <= 23;
        X[55] <= 241;
        out   <= 0;
    end else begin
        X[1]  <= 236;
        X[2]  <= 184;
        X[3]  <= 170;
        X[4]  <= 59;
        X[5]  <= 95;
        X[6]  <= 72;
        X[7]  <= 210;
        X[8]  <= 119;
        X[9]  <= 219;
        X[10] <= 230;
        X[11] <= 74;
        X[12] <= 107;
        X[13] <= 160;
        X[14] <= 44;
        X[15] <= 131;
        X[16] <= 190;
        X[17] <= 246;
        X[18] <= 6;
        X[19] <= 121;
        X[20] <= 76;
        X[21] <= 5;
        X[22] <= 144;
        X[23] <= 193;
        X[24] <= 84;
        X[25] <= 12;
        X[26] <= 255;
        X[27] <= 107;
        X[28] <= 41;
        X[29] <= 43;
        X[30] <= 134;
        X[31] <= 228;
        X[32] <= 134;
        X[33] <= 157;
        X[34] <= 219;
        X[35] <= 106;
        X[36] <= 45;
        X[37] <= 192;
        X[38] <= 142;
        X[39] <= 218;
        X[40] <= 193;
        X[41] <= 173;
        X[42] <= 23;
        X[43] <= 163;
        X[44] <= 63;
        X[45] <= 133;
        X[46] <= 216;
        X[47] <= 60;
        X[48] <= 184;
        X[49] <= 147;
        X[50] <= 129;
        X[51] <= 133;
        X[52] <= 241;
        X[53] <= 63;
        X[54] <= 243;
        X[55] <= 22;
        out   <= 0;
    end
end else begin
    X[55] <= X[54];
    X[54] <= X[53];
    X[53] <= X[52];
    X[52] <= X[51];
    X[51] <= X[50];
    X[50] <= X[49];
    X[49] <= X[48];
    X[48] <= X[47];
    X[47] <= X[46];
    X[46] <= X[45];
    X[45] <= X[44];
    X[44] <= X[43];
    X[43] <= X[42];
    X[42] <= X[41];
    X[41] <= X[40];
    X[40] <= X[39];
    X[39] <= X[38];
    X[38] <= X[37];
    X[37] <= X[36];
    X[36] <= X[35];
    X[35] <= X[34];
    X[34] <= X[33];
    X[33] <= X[32];
    X[32] <= X[31];
    X[31] <= X[30];
    X[30] <= X[29];
    X[29] <= X[28];
    X[28] <= X[27];
    X[27] <= X[26];
    X[26] <= X[25];
    X[25] <= X[24];
    X[24] <= X[23];
    X[23] <= X[22];
    X[22] <= X[21];
    X[21] <= X[20];
    X[20] <= X[19];
    X[19] <= X[18];
    X[18] <= X[17];
    X[17] <= X[16];
    X[16] <= X[15];
    X[15] <= X[14];
    X[14] <= X[13];
    X[13] <= X[12];
    X[12] <= X[11];
    X[11] <= X[10];
    X[10] <= X[9];
    X[9]  <= X[8];
    X[8]  <= X[7];
    X[7]  <= X[6];
    X[6]  <= X[5];
    X[5]  <= X[4];
    X[4]  <= X[3];
    X[3]  <= X[2];
    X[2]  <= X[1];
    X[1]  <= X[55] - X[24];
    out   <= X[1];
end
endgenerate

endmodule
