`ifndef FIR_SYST_SVH
`define FIR_SYST_SVH

`include "macro.svh"
`include "fir.svh"

`define FIR_SYST_ID_CONST  (16'h18DD)

`endif