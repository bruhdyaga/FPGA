module ch_mul_rom(
    input              clk,
    output logic [9:0] data,
    input        [8:0] addr
);

always_ff@(posedge clk) begin
    case (addr)
        {2'b11, 2'b11, 5'd0}      : data <= {-5'd11, -5'd11};
        {2'b11, 2'b11, 5'd1}      : data <= {-5'd12, -5'd8};
        {2'b11, 2'b11, 5'd2}      : data <= {-5'd14, -5'd6};
        {2'b11, 2'b11, 5'd3}      : data <= {-5'd15, -5'd3};
        {2'b11, 2'b11, 5'd4}      : data <= {-5'd15, 5'd0};
        {2'b11, 2'b11, 5'd5}      : data <= {-5'd15, 5'd3};
        {2'b11, 2'b11, 5'd6}      : data <= {-5'd14, 5'd6};
        {2'b11, 2'b11, 5'd7}      : data <= {-5'd12, 5'd8};
        {2'b11, 2'b11, 5'd8}      : data <= {-5'd11, 5'd11};
        {2'b11, 2'b11, 5'd9}      : data <= {-5'd8, 5'd12};
        {2'b11, 2'b11, 5'd10}     : data <= {-5'd6, 5'd14};
        {2'b11, 2'b11, 5'd11}     : data <= {-5'd3, 5'd15};
        {2'b11, 2'b11, 5'd12}     : data <= {5'd0, 5'd15};
        {2'b11, 2'b11, 5'd13}     : data <= {5'd3, 5'd15};
        {2'b11, 2'b11, 5'd14}     : data <= {5'd6, 5'd14};
        {2'b11, 2'b11, 5'd15}     : data <= {5'd8, 5'd12};
        {2'b11, 2'b11, 5'd16}     : data <= {5'd11, 5'd11};
        {2'b11, 2'b11, 5'd17}     : data <= {5'd12, 5'd8};
        {2'b11, 2'b11, 5'd18}     : data <= {5'd14, 5'd6};
        {2'b11, 2'b11, 5'd19}     : data <= {5'd15, 5'd3};
        {2'b11, 2'b11, 5'd20}     : data <= {5'd15, 5'd0};
        {2'b11, 2'b11, 5'd21}     : data <= {5'd15, -5'd3};
        {2'b11, 2'b11, 5'd22}     : data <= {5'd14, -5'd6};
        {2'b11, 2'b11, 5'd23}     : data <= {5'd12, -5'd8};
        {2'b11, 2'b11, 5'd24}     : data <= {5'd11, -5'd11};
        {2'b11, 2'b11, 5'd25}     : data <= {5'd8, -5'd12};
        {2'b11, 2'b11, 5'd26}     : data <= {5'd6, -5'd14};
        {2'b11, 2'b11, 5'd27}     : data <= {5'd3, -5'd15};
        {2'b11, 2'b11, 5'd28}     : data <= {5'd0, -5'd15};
        {2'b11, 2'b11, 5'd29}     : data <= {-5'd3, -5'd15};
        {2'b11, 2'b11, 5'd30}     : data <= {-5'd6, -5'd14};
        {2'b11, 2'b11, 5'd31}     : data <= {-5'd8, -5'd12};
        
        {2'b11, 2'b10, 5'd0}      : data <= {-5'd11, -5'd4};
        {2'b11, 2'b10, 5'd1}      : data <= {-5'd11, -5'd1};
        {2'b11, 2'b10, 5'd2}      : data <= {-5'd11, 5'd1};
        {2'b11, 2'b10, 5'd3}      : data <= {-5'd11, 5'd3};
        {2'b11, 2'b10, 5'd4}      : data <= {-5'd10, 5'd5};
        {2'b11, 2'b10, 5'd5}      : data <= {-5'd9, 5'd7};
        {2'b11, 2'b10, 5'd6}      : data <= {-5'd7, 5'd8};
        {2'b11, 2'b10, 5'd7}      : data <= {-5'd6, 5'd10};
        {2'b11, 2'b10, 5'd8}      : data <= {-5'd4, 5'd11};
        {2'b11, 2'b10, 5'd9}      : data <= {-5'd1, 5'd11};
        {2'b11, 2'b10, 5'd10}     : data <= {5'd1, 5'd11};
        {2'b11, 2'b10, 5'd11}     : data <= {5'd3, 5'd11};
        {2'b11, 2'b10, 5'd12}     : data <= {5'd5, 5'd10};
        {2'b11, 2'b10, 5'd13}     : data <= {5'd7, 5'd9};
        {2'b11, 2'b10, 5'd14}     : data <= {5'd8, 5'd7};
        {2'b11, 2'b10, 5'd15}     : data <= {5'd10, 5'd6};
        {2'b11, 2'b10, 5'd16}     : data <= {5'd11, 5'd4};
        {2'b11, 2'b10, 5'd17}     : data <= {5'd11, 5'd1};
        {2'b11, 2'b10, 5'd18}     : data <= {5'd11, -5'd1};
        {2'b11, 2'b10, 5'd19}     : data <= {5'd11, -5'd3};
        {2'b11, 2'b10, 5'd20}     : data <= {5'd10, -5'd5};
        {2'b11, 2'b10, 5'd21}     : data <= {5'd9, -5'd7};
        {2'b11, 2'b10, 5'd22}     : data <= {5'd7, -5'd8};
        {2'b11, 2'b10, 5'd23}     : data <= {5'd6, -5'd10};
        {2'b11, 2'b10, 5'd24}     : data <= {5'd4, -5'd11};
        {2'b11, 2'b10, 5'd25}     : data <= {5'd1, -5'd11};
        {2'b11, 2'b10, 5'd26}     : data <= {-5'd1, -5'd11};
        {2'b11, 2'b10, 5'd27}     : data <= {-5'd3, -5'd11};
        {2'b11, 2'b10, 5'd28}     : data <= {-5'd5, -5'd10};
        {2'b11, 2'b10, 5'd29}     : data <= {-5'd7, -5'd9};
        {2'b11, 2'b10, 5'd30}     : data <= {-5'd8, -5'd7};
        {2'b11, 2'b10, 5'd31}     : data <= {-5'd10, -5'd6};
        
        {2'b11, 2'b00, 5'd0}      : data <= {-5'd11, 5'd4};
        {2'b11, 2'b00, 5'd1}      : data <= {-5'd10, 5'd6};
        {2'b11, 2'b00, 5'd2}      : data <= {-5'd8, 5'd7};
        {2'b11, 2'b00, 5'd3}      : data <= {-5'd7, 5'd9};
        {2'b11, 2'b00, 5'd4}      : data <= {-5'd5, 5'd10};
        {2'b11, 2'b00, 5'd5}      : data <= {-5'd3, 5'd11};
        {2'b11, 2'b00, 5'd6}      : data <= {-5'd1, 5'd11};
        {2'b11, 2'b00, 5'd7}      : data <= {5'd1, 5'd11};
        {2'b11, 2'b00, 5'd8}      : data <= {5'd4, 5'd11};
        {2'b11, 2'b00, 5'd9}      : data <= {5'd6, 5'd10};
        {2'b11, 2'b00, 5'd10}     : data <= {5'd7, 5'd8};
        {2'b11, 2'b00, 5'd11}     : data <= {5'd9, 5'd7};
        {2'b11, 2'b00, 5'd12}     : data <= {5'd10, 5'd5};
        {2'b11, 2'b00, 5'd13}     : data <= {5'd11, 5'd3};
        {2'b11, 2'b00, 5'd14}     : data <= {5'd11, 5'd1};
        {2'b11, 2'b00, 5'd15}     : data <= {5'd11, -5'd1};
        {2'b11, 2'b00, 5'd16}     : data <= {5'd11, -5'd4};
        {2'b11, 2'b00, 5'd17}     : data <= {5'd10, -5'd6};
        {2'b11, 2'b00, 5'd18}     : data <= {5'd8, -5'd7};
        {2'b11, 2'b00, 5'd19}     : data <= {5'd7, -5'd9};
        {2'b11, 2'b00, 5'd20}     : data <= {5'd5, -5'd10};
        {2'b11, 2'b00, 5'd21}     : data <= {5'd3, -5'd11};
        {2'b11, 2'b00, 5'd22}     : data <= {5'd1, -5'd11};
        {2'b11, 2'b00, 5'd23}     : data <= {-5'd1, -5'd11};
        {2'b11, 2'b00, 5'd24}     : data <= {-5'd4, -5'd11};
        {2'b11, 2'b00, 5'd25}     : data <= {-5'd6, -5'd10};
        {2'b11, 2'b00, 5'd26}     : data <= {-5'd7, -5'd8};
        {2'b11, 2'b00, 5'd27}     : data <= {-5'd9, -5'd7};
        {2'b11, 2'b00, 5'd28}     : data <= {-5'd10, -5'd5};
        {2'b11, 2'b00, 5'd29}     : data <= {-5'd11, -5'd3};
        {2'b11, 2'b00, 5'd30}     : data <= {-5'd11, -5'd1};
        {2'b11, 2'b00, 5'd31}     : data <= {-5'd11, 5'd1};
        
        {2'b11, 2'b01, 5'd0}      : data <= {-5'd11, 5'd11};
        {2'b11, 2'b01, 5'd1}      : data <= {-5'd8, 5'd12};
        {2'b11, 2'b01, 5'd2}      : data <= {-5'd6, 5'd14};
        {2'b11, 2'b01, 5'd3}      : data <= {-5'd3, 5'd15};
        {2'b11, 2'b01, 5'd4}      : data <= {5'd0, 5'd15};
        {2'b11, 2'b01, 5'd5}      : data <= {5'd3, 5'd15};
        {2'b11, 2'b01, 5'd6}      : data <= {5'd6, 5'd14};
        {2'b11, 2'b01, 5'd7}      : data <= {5'd8, 5'd12};
        {2'b11, 2'b01, 5'd8}      : data <= {5'd11, 5'd11};
        {2'b11, 2'b01, 5'd9}      : data <= {5'd12, 5'd8};
        {2'b11, 2'b01, 5'd10}     : data <= {5'd14, 5'd6};
        {2'b11, 2'b01, 5'd11}     : data <= {5'd15, 5'd3};
        {2'b11, 2'b01, 5'd12}     : data <= {5'd15, 5'd0};
        {2'b11, 2'b01, 5'd13}     : data <= {5'd15, -5'd3};
        {2'b11, 2'b01, 5'd14}     : data <= {5'd14, -5'd6};
        {2'b11, 2'b01, 5'd15}     : data <= {5'd12, -5'd8};
        {2'b11, 2'b01, 5'd16}     : data <= {5'd11, -5'd11};
        {2'b11, 2'b01, 5'd17}     : data <= {5'd8, -5'd12};
        {2'b11, 2'b01, 5'd18}     : data <= {5'd6, -5'd14};
        {2'b11, 2'b01, 5'd19}     : data <= {5'd3, -5'd15};
        {2'b11, 2'b01, 5'd20}     : data <= {5'd0, -5'd15};
        {2'b11, 2'b01, 5'd21}     : data <= {-5'd3, -5'd15};
        {2'b11, 2'b01, 5'd22}     : data <= {-5'd6, -5'd14};
        {2'b11, 2'b01, 5'd23}     : data <= {-5'd8, -5'd12};
        {2'b11, 2'b01, 5'd24}     : data <= {-5'd11, -5'd11};
        {2'b11, 2'b01, 5'd25}     : data <= {-5'd12, -5'd8};
        {2'b11, 2'b01, 5'd26}     : data <= {-5'd14, -5'd6};
        {2'b11, 2'b01, 5'd27}     : data <= {-5'd15, -5'd3};
        {2'b11, 2'b01, 5'd28}     : data <= {-5'd15, 5'd0};
        {2'b11, 2'b01, 5'd29}     : data <= {-5'd15, 5'd3};
        {2'b11, 2'b01, 5'd30}     : data <= {-5'd14, 5'd6};
        {2'b11, 2'b01, 5'd31}     : data <= {-5'd12, 5'd8};
        
        
        {2'b10, 2'b11, 5'd0}      : data <= {-5'd4, -5'd11};
        {2'b10, 2'b11, 5'd1}      : data <= {-5'd6, -5'd10};
        {2'b10, 2'b11, 5'd2}      : data <= {-5'd7, -5'd8};
        {2'b10, 2'b11, 5'd3}      : data <= {-5'd9, -5'd7};
        {2'b10, 2'b11, 5'd4}      : data <= {-5'd10, -5'd5};
        {2'b10, 2'b11, 5'd5}      : data <= {-5'd11, -5'd3};
        {2'b10, 2'b11, 5'd6}      : data <= {-5'd11, -5'd1};
        {2'b10, 2'b11, 5'd7}      : data <= {-5'd11, 5'd1};
        {2'b10, 2'b11, 5'd8}      : data <= {-5'd11, 5'd4};
        {2'b10, 2'b11, 5'd9}      : data <= {-5'd10, 5'd6};
        {2'b10, 2'b11, 5'd10}     : data <= {-5'd8, 5'd7};
        {2'b10, 2'b11, 5'd11}     : data <= {-5'd7, 5'd9};
        {2'b10, 2'b11, 5'd12}     : data <= {-5'd5, 5'd10};
        {2'b10, 2'b11, 5'd13}     : data <= {-5'd3, 5'd11};
        {2'b10, 2'b11, 5'd14}     : data <= {-5'd1, 5'd11};
        {2'b10, 2'b11, 5'd15}     : data <= {5'd1, 5'd11};
        {2'b10, 2'b11, 5'd16}     : data <= {5'd4, 5'd11};
        {2'b10, 2'b11, 5'd17}     : data <= {5'd6, 5'd10};
        {2'b10, 2'b11, 5'd18}     : data <= {5'd7, 5'd8};
        {2'b10, 2'b11, 5'd19}     : data <= {5'd9, 5'd7};
        {2'b10, 2'b11, 5'd20}     : data <= {5'd10, 5'd5};
        {2'b10, 2'b11, 5'd21}     : data <= {5'd11, 5'd3};
        {2'b10, 2'b11, 5'd22}     : data <= {5'd11, 5'd1};
        {2'b10, 2'b11, 5'd23}     : data <= {5'd11, -5'd1};
        {2'b10, 2'b11, 5'd24}     : data <= {5'd11, -5'd4};
        {2'b10, 2'b11, 5'd25}     : data <= {5'd10, -5'd6};
        {2'b10, 2'b11, 5'd26}     : data <= {5'd8, -5'd7};
        {2'b10, 2'b11, 5'd27}     : data <= {5'd7, -5'd9};
        {2'b10, 2'b11, 5'd28}     : data <= {5'd5, -5'd10};
        {2'b10, 2'b11, 5'd29}     : data <= {5'd3, -5'd11};
        {2'b10, 2'b11, 5'd30}     : data <= {5'd1, -5'd11};
        {2'b10, 2'b11, 5'd31}     : data <= {-5'd1, -5'd11};
        
        {2'b10, 2'b10, 5'd0}      : data <= {-5'd4, -5'd4};
        {2'b10, 2'b10, 5'd1}      : data <= {-5'd4, -5'd3};
        {2'b10, 2'b10, 5'd2}      : data <= {-5'd5, -5'd2};
        {2'b10, 2'b10, 5'd3}      : data <= {-5'd5, -5'd1};
        {2'b10, 2'b10, 5'd4}      : data <= {-5'd5, 5'd0};
        {2'b10, 2'b10, 5'd5}      : data <= {-5'd5, 5'd1};
        {2'b10, 2'b10, 5'd6}      : data <= {-5'd5, 5'd2};
        {2'b10, 2'b10, 5'd7}      : data <= {-5'd4, 5'd3};
        {2'b10, 2'b10, 5'd8}      : data <= {-5'd4, 5'd4};
        {2'b10, 2'b10, 5'd9}      : data <= {-5'd3, 5'd4};
        {2'b10, 2'b10, 5'd10}     : data <= {-5'd2, 5'd5};
        {2'b10, 2'b10, 5'd11}     : data <= {-5'd1, 5'd5};
        {2'b10, 2'b10, 5'd12}     : data <= {5'd0, 5'd5};
        {2'b10, 2'b10, 5'd13}     : data <= {5'd1, 5'd5};
        {2'b10, 2'b10, 5'd14}     : data <= {5'd2, 5'd5};
        {2'b10, 2'b10, 5'd15}     : data <= {5'd3, 5'd4};
        {2'b10, 2'b10, 5'd16}     : data <= {5'd4, 5'd4};
        {2'b10, 2'b10, 5'd17}     : data <= {5'd4, 5'd3};
        {2'b10, 2'b10, 5'd18}     : data <= {5'd5, 5'd2};
        {2'b10, 2'b10, 5'd19}     : data <= {5'd5, 5'd1};
        {2'b10, 2'b10, 5'd20}     : data <= {5'd5, 5'd0};
        {2'b10, 2'b10, 5'd21}     : data <= {5'd5, -5'd1};
        {2'b10, 2'b10, 5'd22}     : data <= {5'd5, -5'd2};
        {2'b10, 2'b10, 5'd23}     : data <= {5'd4, -5'd3};
        {2'b10, 2'b10, 5'd24}     : data <= {5'd4, -5'd4};
        {2'b10, 2'b10, 5'd25}     : data <= {5'd3, -5'd4};
        {2'b10, 2'b10, 5'd26}     : data <= {5'd2, -5'd5};
        {2'b10, 2'b10, 5'd27}     : data <= {5'd1, -5'd5};
        {2'b10, 2'b10, 5'd28}     : data <= {5'd0, -5'd5};
        {2'b10, 2'b10, 5'd29}     : data <= {-5'd1, -5'd5};
        {2'b10, 2'b10, 5'd30}     : data <= {-5'd2, -5'd5};
        {2'b10, 2'b10, 5'd31}     : data <= {-5'd3, -5'd4};
        
        {2'b10, 2'b00, 5'd0}      : data <= {-5'd4, 5'd4};
        {2'b10, 2'b00, 5'd1}      : data <= {-5'd3, 5'd4};
        {2'b10, 2'b00, 5'd2}      : data <= {-5'd2, 5'd5};
        {2'b10, 2'b00, 5'd3}      : data <= {-5'd1, 5'd5};
        {2'b10, 2'b00, 5'd4}      : data <= {5'd0, 5'd5};
        {2'b10, 2'b00, 5'd5}      : data <= {5'd1, 5'd5};
        {2'b10, 2'b00, 5'd6}      : data <= {5'd2, 5'd5};
        {2'b10, 2'b00, 5'd7}      : data <= {5'd3, 5'd4};
        {2'b10, 2'b00, 5'd8}      : data <= {5'd4, 5'd4};
        {2'b10, 2'b00, 5'd9}      : data <= {5'd4, 5'd3};
        {2'b10, 2'b00, 5'd10}     : data <= {5'd5, 5'd2};
        {2'b10, 2'b00, 5'd11}     : data <= {5'd5, 5'd1};
        {2'b10, 2'b00, 5'd12}     : data <= {5'd5, 5'd0};
        {2'b10, 2'b00, 5'd13}     : data <= {5'd5, -5'd1};
        {2'b10, 2'b00, 5'd14}     : data <= {5'd5, -5'd2};
        {2'b10, 2'b00, 5'd15}     : data <= {5'd4, -5'd3};
        {2'b10, 2'b00, 5'd16}     : data <= {5'd4, -5'd4};
        {2'b10, 2'b00, 5'd17}     : data <= {5'd3, -5'd4};
        {2'b10, 2'b00, 5'd18}     : data <= {5'd2, -5'd5};
        {2'b10, 2'b00, 5'd19}     : data <= {5'd1, -5'd5};
        {2'b10, 2'b00, 5'd20}     : data <= {5'd0, -5'd5};
        {2'b10, 2'b00, 5'd21}     : data <= {-5'd1, -5'd5};
        {2'b10, 2'b00, 5'd22}     : data <= {-5'd2, -5'd5};
        {2'b10, 2'b00, 5'd23}     : data <= {-5'd3, -5'd4};
        {2'b10, 2'b00, 5'd24}     : data <= {-5'd4, -5'd4};
        {2'b10, 2'b00, 5'd25}     : data <= {-5'd4, -5'd3};
        {2'b10, 2'b00, 5'd26}     : data <= {-5'd5, -5'd2};
        {2'b10, 2'b00, 5'd27}     : data <= {-5'd5, -5'd1};
        {2'b10, 2'b00, 5'd28}     : data <= {-5'd5, 5'd0};
        {2'b10, 2'b00, 5'd29}     : data <= {-5'd5, 5'd1};
        {2'b10, 2'b00, 5'd30}     : data <= {-5'd5, 5'd2};
        {2'b10, 2'b00, 5'd31}     : data <= {-5'd4, 5'd3};
        
        {2'b10, 2'b01, 5'd0}      : data <= {-5'd4, 5'd11};
        {2'b10, 2'b01, 5'd1}      : data <= {-5'd1, 5'd11};
        {2'b10, 2'b01, 5'd2}      : data <= {5'd1, 5'd11};
        {2'b10, 2'b01, 5'd3}      : data <= {5'd3, 5'd11};
        {2'b10, 2'b01, 5'd4}      : data <= {5'd5, 5'd10};
        {2'b10, 2'b01, 5'd5}      : data <= {5'd7, 5'd9};
        {2'b10, 2'b01, 5'd6}      : data <= {5'd8, 5'd7};
        {2'b10, 2'b01, 5'd7}      : data <= {5'd10, 5'd6};
        {2'b10, 2'b01, 5'd8}      : data <= {5'd11, 5'd4};
        {2'b10, 2'b01, 5'd9}      : data <= {5'd11, 5'd1};
        {2'b10, 2'b01, 5'd10}     : data <= {5'd11, -5'd1};
        {2'b10, 2'b01, 5'd11}     : data <= {5'd11, -5'd3};
        {2'b10, 2'b01, 5'd12}     : data <= {5'd10, -5'd5};
        {2'b10, 2'b01, 5'd13}     : data <= {5'd9, -5'd7};
        {2'b10, 2'b01, 5'd14}     : data <= {5'd7, -5'd8};
        {2'b10, 2'b01, 5'd15}     : data <= {5'd6, -5'd10};
        {2'b10, 2'b01, 5'd16}     : data <= {5'd4, -5'd11};
        {2'b10, 2'b01, 5'd17}     : data <= {5'd1, -5'd11};
        {2'b10, 2'b01, 5'd18}     : data <= {-5'd1, -5'd11};
        {2'b10, 2'b01, 5'd19}     : data <= {-5'd3, -5'd11};
        {2'b10, 2'b01, 5'd20}     : data <= {-5'd5, -5'd10};
        {2'b10, 2'b01, 5'd21}     : data <= {-5'd7, -5'd9};
        {2'b10, 2'b01, 5'd22}     : data <= {-5'd8, -5'd7};
        {2'b10, 2'b01, 5'd23}     : data <= {-5'd10, -5'd6};
        {2'b10, 2'b01, 5'd24}     : data <= {-5'd11, -5'd4};
        {2'b10, 2'b01, 5'd25}     : data <= {-5'd11, -5'd1};
        {2'b10, 2'b01, 5'd26}     : data <= {-5'd11, 5'd1};
        {2'b10, 2'b01, 5'd27}     : data <= {-5'd11, 5'd3};
        {2'b10, 2'b01, 5'd28}     : data <= {-5'd10, 5'd5};
        {2'b10, 2'b01, 5'd29}     : data <= {-5'd9, 5'd7};
        {2'b10, 2'b01, 5'd30}     : data <= {-5'd7, 5'd8};
        {2'b10, 2'b01, 5'd31}     : data <= {-5'd6, 5'd10};
        
        
        {2'b00, 2'b11, 5'd0}      : data <= {5'd4, -5'd11};
        {2'b00, 2'b11, 5'd1}      : data <= {5'd1, -5'd11};
        {2'b00, 2'b11, 5'd2}      : data <= {-5'd1, -5'd11};
        {2'b00, 2'b11, 5'd3}      : data <= {-5'd3, -5'd11};
        {2'b00, 2'b11, 5'd4}      : data <= {-5'd5, -5'd10};
        {2'b00, 2'b11, 5'd5}      : data <= {-5'd7, -5'd9};
        {2'b00, 2'b11, 5'd6}      : data <= {-5'd8, -5'd7};
        {2'b00, 2'b11, 5'd7}      : data <= {-5'd10, -5'd6};
        {2'b00, 2'b11, 5'd8}      : data <= {-5'd11, -5'd4};
        {2'b00, 2'b11, 5'd9}      : data <= {-5'd11, -5'd1};
        {2'b00, 2'b11, 5'd10}     : data <= {-5'd11, 5'd1};
        {2'b00, 2'b11, 5'd11}     : data <= {-5'd11, 5'd3};
        {2'b00, 2'b11, 5'd12}     : data <= {-5'd10, 5'd5};
        {2'b00, 2'b11, 5'd13}     : data <= {-5'd9, 5'd7};
        {2'b00, 2'b11, 5'd14}     : data <= {-5'd7, 5'd8};
        {2'b00, 2'b11, 5'd15}     : data <= {-5'd6, 5'd10};
        {2'b00, 2'b11, 5'd16}     : data <= {-5'd4, 5'd11};
        {2'b00, 2'b11, 5'd17}     : data <= {-5'd1, 5'd11};
        {2'b00, 2'b11, 5'd18}     : data <= {5'd1, 5'd11};
        {2'b00, 2'b11, 5'd19}     : data <= {5'd3, 5'd11};
        {2'b00, 2'b11, 5'd20}     : data <= {5'd5, 5'd10};
        {2'b00, 2'b11, 5'd21}     : data <= {5'd7, 5'd9};
        {2'b00, 2'b11, 5'd22}     : data <= {5'd8, 5'd7};
        {2'b00, 2'b11, 5'd23}     : data <= {5'd10, 5'd6};
        {2'b00, 2'b11, 5'd24}     : data <= {5'd11, 5'd4};
        {2'b00, 2'b11, 5'd25}     : data <= {5'd11, 5'd1};
        {2'b00, 2'b11, 5'd26}     : data <= {5'd11, -5'd1};
        {2'b00, 2'b11, 5'd27}     : data <= {5'd11, -5'd3};
        {2'b00, 2'b11, 5'd28}     : data <= {5'd10, -5'd5};
        {2'b00, 2'b11, 5'd29}     : data <= {5'd9, -5'd7};
        {2'b00, 2'b11, 5'd30}     : data <= {5'd7, -5'd8};
        {2'b00, 2'b11, 5'd31}     : data <= {5'd6, -5'd10};
        
        {2'b00, 2'b10, 5'd0}      : data <= {5'd4, -5'd4};
        {2'b00, 2'b10, 5'd1}      : data <= {5'd3, -5'd4};
        {2'b00, 2'b10, 5'd2}      : data <= {5'd2, -5'd5};
        {2'b00, 2'b10, 5'd3}      : data <= {5'd1, -5'd5};
        {2'b00, 2'b10, 5'd4}      : data <= {5'd0, -5'd5};
        {2'b00, 2'b10, 5'd5}      : data <= {-5'd1, -5'd5};
        {2'b00, 2'b10, 5'd6}      : data <= {-5'd2, -5'd5};
        {2'b00, 2'b10, 5'd7}      : data <= {-5'd3, -5'd4};
        {2'b00, 2'b10, 5'd8}      : data <= {-5'd4, -5'd4};
        {2'b00, 2'b10, 5'd9}      : data <= {-5'd4, -5'd3};
        {2'b00, 2'b10, 5'd10}     : data <= {-5'd5, -5'd2};
        {2'b00, 2'b10, 5'd11}     : data <= {-5'd5, -5'd1};
        {2'b00, 2'b10, 5'd12}     : data <= {-5'd5, 5'd0};
        {2'b00, 2'b10, 5'd13}     : data <= {-5'd5, 5'd1};
        {2'b00, 2'b10, 5'd14}     : data <= {-5'd5, 5'd2};
        {2'b00, 2'b10, 5'd15}     : data <= {-5'd4, 5'd3};
        {2'b00, 2'b10, 5'd16}     : data <= {-5'd4, 5'd4};
        {2'b00, 2'b10, 5'd17}     : data <= {-5'd3, 5'd4};
        {2'b00, 2'b10, 5'd18}     : data <= {-5'd2, 5'd5};
        {2'b00, 2'b10, 5'd19}     : data <= {-5'd1, 5'd5};
        {2'b00, 2'b10, 5'd20}     : data <= {5'd0, 5'd5};
        {2'b00, 2'b10, 5'd21}     : data <= {5'd1, 5'd5};
        {2'b00, 2'b10, 5'd22}     : data <= {5'd2, 5'd5};
        {2'b00, 2'b10, 5'd23}     : data <= {5'd3, 5'd4};
        {2'b00, 2'b10, 5'd24}     : data <= {5'd4, 5'd4};
        {2'b00, 2'b10, 5'd25}     : data <= {5'd4, 5'd3};
        {2'b00, 2'b10, 5'd26}     : data <= {5'd5, 5'd2};
        {2'b00, 2'b10, 5'd27}     : data <= {5'd5, 5'd1};
        {2'b00, 2'b10, 5'd28}     : data <= {5'd5, 5'd0};
        {2'b00, 2'b10, 5'd29}     : data <= {5'd5, -5'd1};
        {2'b00, 2'b10, 5'd30}     : data <= {5'd5, -5'd2};
        {2'b00, 2'b10, 5'd31}     : data <= {5'd4, -5'd3};
        
        {2'b00, 2'b00, 5'd0}      : data <= {5'd4, 5'd4};
        {2'b00, 2'b00, 5'd1}      : data <= {5'd4, 5'd3};
        {2'b00, 2'b00, 5'd2}      : data <= {5'd5, 5'd2};
        {2'b00, 2'b00, 5'd3}      : data <= {5'd5, 5'd1};
        {2'b00, 2'b00, 5'd4}      : data <= {5'd5, 5'd0};
        {2'b00, 2'b00, 5'd5}      : data <= {5'd5, -5'd1};
        {2'b00, 2'b00, 5'd6}      : data <= {5'd5, -5'd2};
        {2'b00, 2'b00, 5'd7}      : data <= {5'd4, -5'd3};
        {2'b00, 2'b00, 5'd8}      : data <= {5'd4, -5'd4};
        {2'b00, 2'b00, 5'd9}      : data <= {5'd3, -5'd4};
        {2'b00, 2'b00, 5'd10}     : data <= {5'd2, -5'd5};
        {2'b00, 2'b00, 5'd11}     : data <= {5'd1, -5'd5};
        {2'b00, 2'b00, 5'd12}     : data <= {5'd0, -5'd5};
        {2'b00, 2'b00, 5'd13}     : data <= {-5'd1, -5'd5};
        {2'b00, 2'b00, 5'd14}     : data <= {-5'd2, -5'd5};
        {2'b00, 2'b00, 5'd15}     : data <= {-5'd3, -5'd4};
        {2'b00, 2'b00, 5'd16}     : data <= {-5'd4, -5'd4};
        {2'b00, 2'b00, 5'd17}     : data <= {-5'd4, -5'd3};
        {2'b00, 2'b00, 5'd18}     : data <= {-5'd5, -5'd2};
        {2'b00, 2'b00, 5'd19}     : data <= {-5'd5, -5'd1};
        {2'b00, 2'b00, 5'd20}     : data <= {-5'd5, 5'd0};
        {2'b00, 2'b00, 5'd21}     : data <= {-5'd5, 5'd1};
        {2'b00, 2'b00, 5'd22}     : data <= {-5'd5, 5'd2};
        {2'b00, 2'b00, 5'd23}     : data <= {-5'd4, 5'd3};
        {2'b00, 2'b00, 5'd24}     : data <= {-5'd4, 5'd4};
        {2'b00, 2'b00, 5'd25}     : data <= {-5'd3, 5'd4};
        {2'b00, 2'b00, 5'd26}     : data <= {-5'd2, 5'd5};
        {2'b00, 2'b00, 5'd27}     : data <= {-5'd1, 5'd5};
        {2'b00, 2'b00, 5'd28}     : data <= {5'd0, 5'd5};
        {2'b00, 2'b00, 5'd29}     : data <= {5'd1, 5'd5};
        {2'b00, 2'b00, 5'd30}     : data <= {5'd2, 5'd5};
        {2'b00, 2'b00, 5'd31}     : data <= {5'd3, 5'd4};
        
        {2'b00, 2'b01, 5'd0}      : data <= {5'd4, 5'd11};
        {2'b00, 2'b01, 5'd1}      : data <= {5'd6, 5'd10};
        {2'b00, 2'b01, 5'd2}      : data <= {5'd7, 5'd8};
        {2'b00, 2'b01, 5'd3}      : data <= {5'd9, 5'd7};
        {2'b00, 2'b01, 5'd4}      : data <= {5'd10, 5'd5};
        {2'b00, 2'b01, 5'd5}      : data <= {5'd11, 5'd3};
        {2'b00, 2'b01, 5'd6}      : data <= {5'd11, 5'd1};
        {2'b00, 2'b01, 5'd7}      : data <= {5'd11, -5'd1};
        {2'b00, 2'b01, 5'd8}      : data <= {5'd11, -5'd4};
        {2'b00, 2'b01, 5'd9}      : data <= {5'd10, -5'd6};
        {2'b00, 2'b01, 5'd10}     : data <= {5'd8, -5'd7};
        {2'b00, 2'b01, 5'd11}     : data <= {5'd7, -5'd9};
        {2'b00, 2'b01, 5'd12}     : data <= {5'd5, -5'd10};
        {2'b00, 2'b01, 5'd13}     : data <= {5'd3, -5'd11};
        {2'b00, 2'b01, 5'd14}     : data <= {5'd1, -5'd11};
        {2'b00, 2'b01, 5'd15}     : data <= {-5'd1, -5'd11};
        {2'b00, 2'b01, 5'd16}     : data <= {-5'd4, -5'd11};
        {2'b00, 2'b01, 5'd17}     : data <= {-5'd6, -5'd10};
        {2'b00, 2'b01, 5'd18}     : data <= {-5'd7, -5'd8};
        {2'b00, 2'b01, 5'd19}     : data <= {-5'd9, -5'd7};
        {2'b00, 2'b01, 5'd20}     : data <= {-5'd10, -5'd5};
        {2'b00, 2'b01, 5'd21}     : data <= {-5'd11, -5'd3};
        {2'b00, 2'b01, 5'd22}     : data <= {-5'd11, -5'd1};
        {2'b00, 2'b01, 5'd23}     : data <= {-5'd11, 5'd1};
        {2'b00, 2'b01, 5'd24}     : data <= {-5'd11, 5'd4};
        {2'b00, 2'b01, 5'd25}     : data <= {-5'd10, 5'd6};
        {2'b00, 2'b01, 5'd26}     : data <= {-5'd8, 5'd7};
        {2'b00, 2'b01, 5'd27}     : data <= {-5'd7, 5'd9};
        {2'b00, 2'b01, 5'd28}     : data <= {-5'd5, 5'd10};
        {2'b00, 2'b01, 5'd29}     : data <= {-5'd3, 5'd11};
        {2'b00, 2'b01, 5'd30}     : data <= {-5'd1, 5'd11};
        {2'b00, 2'b01, 5'd31}     : data <= {5'd1, 5'd11};
        
        
        {2'b01, 2'b11, 5'd0}      : data <= {5'd11, -5'd11};
        {2'b01, 2'b11, 5'd1}      : data <= {5'd8, -5'd12};
        {2'b01, 2'b11, 5'd2}      : data <= {5'd6, -5'd14};
        {2'b01, 2'b11, 5'd3}      : data <= {5'd3, -5'd15};
        {2'b01, 2'b11, 5'd4}      : data <= {5'd0, -5'd15};
        {2'b01, 2'b11, 5'd5}      : data <= {-5'd3, -5'd15};
        {2'b01, 2'b11, 5'd6}      : data <= {-5'd6, -5'd14};
        {2'b01, 2'b11, 5'd7}      : data <= {-5'd8, -5'd12};
        {2'b01, 2'b11, 5'd8}      : data <= {-5'd11, -5'd11};
        {2'b01, 2'b11, 5'd9}      : data <= {-5'd12, -5'd8};
        {2'b01, 2'b11, 5'd10}     : data <= {-5'd14, -5'd6};
        {2'b01, 2'b11, 5'd11}     : data <= {-5'd15, -5'd3};
        {2'b01, 2'b11, 5'd12}     : data <= {-5'd15, 5'd0};
        {2'b01, 2'b11, 5'd13}     : data <= {-5'd15, 5'd3};
        {2'b01, 2'b11, 5'd14}     : data <= {-5'd14, 5'd6};
        {2'b01, 2'b11, 5'd15}     : data <= {-5'd12, 5'd8};
        {2'b01, 2'b11, 5'd16}     : data <= {-5'd11, 5'd11};
        {2'b01, 2'b11, 5'd17}     : data <= {-5'd8, 5'd12};
        {2'b01, 2'b11, 5'd18}     : data <= {-5'd6, 5'd14};
        {2'b01, 2'b11, 5'd19}     : data <= {-5'd3, 5'd15};
        {2'b01, 2'b11, 5'd20}     : data <= {5'd0, 5'd15};
        {2'b01, 2'b11, 5'd21}     : data <= {5'd3, 5'd15};
        {2'b01, 2'b11, 5'd22}     : data <= {5'd6, 5'd14};
        {2'b01, 2'b11, 5'd23}     : data <= {5'd8, 5'd12};
        {2'b01, 2'b11, 5'd24}     : data <= {5'd11, 5'd11};
        {2'b01, 2'b11, 5'd25}     : data <= {5'd12, 5'd8};
        {2'b01, 2'b11, 5'd26}     : data <= {5'd14, 5'd6};
        {2'b01, 2'b11, 5'd27}     : data <= {5'd15, 5'd3};
        {2'b01, 2'b11, 5'd28}     : data <= {5'd15, 5'd0};
        {2'b01, 2'b11, 5'd29}     : data <= {5'd15, -5'd3};
        {2'b01, 2'b11, 5'd30}     : data <= {5'd14, -5'd6};
        {2'b01, 2'b11, 5'd31}     : data <= {5'd12, -5'd8};
        
        {2'b01, 2'b10, 5'd0}      : data <= {5'd11, -5'd4};
        {2'b01, 2'b10, 5'd1}      : data <= {5'd10, -5'd6};
        {2'b01, 2'b10, 5'd2}      : data <= {5'd8, -5'd7};
        {2'b01, 2'b10, 5'd3}      : data <= {5'd7, -5'd9};
        {2'b01, 2'b10, 5'd4}      : data <= {5'd5, -5'd10};
        {2'b01, 2'b10, 5'd5}      : data <= {5'd3, -5'd11};
        {2'b01, 2'b10, 5'd6}      : data <= {5'd1, -5'd11};
        {2'b01, 2'b10, 5'd7}      : data <= {-5'd1, -5'd11};
        {2'b01, 2'b10, 5'd8}      : data <= {-5'd4, -5'd11};
        {2'b01, 2'b10, 5'd9}      : data <= {-5'd6, -5'd10};
        {2'b01, 2'b10, 5'd10}     : data <= {-5'd7, -5'd8};
        {2'b01, 2'b10, 5'd11}     : data <= {-5'd9, -5'd7};
        {2'b01, 2'b10, 5'd12}     : data <= {-5'd10, -5'd5};
        {2'b01, 2'b10, 5'd13}     : data <= {-5'd11, -5'd3};
        {2'b01, 2'b10, 5'd14}     : data <= {-5'd11, -5'd1};
        {2'b01, 2'b10, 5'd15}     : data <= {-5'd11, 5'd1};
        {2'b01, 2'b10, 5'd16}     : data <= {-5'd11, 5'd4};
        {2'b01, 2'b10, 5'd17}     : data <= {-5'd10, 5'd6};
        {2'b01, 2'b10, 5'd18}     : data <= {-5'd8, 5'd7};
        {2'b01, 2'b10, 5'd19}     : data <= {-5'd7, 5'd9};
        {2'b01, 2'b10, 5'd20}     : data <= {-5'd5, 5'd10};
        {2'b01, 2'b10, 5'd21}     : data <= {-5'd3, 5'd11};
        {2'b01, 2'b10, 5'd22}     : data <= {-5'd1, 5'd11};
        {2'b01, 2'b10, 5'd23}     : data <= {5'd1, 5'd11};
        {2'b01, 2'b10, 5'd24}     : data <= {5'd4, 5'd11};
        {2'b01, 2'b10, 5'd25}     : data <= {5'd6, 5'd10};
        {2'b01, 2'b10, 5'd26}     : data <= {5'd7, 5'd8};
        {2'b01, 2'b10, 5'd27}     : data <= {5'd9, 5'd7};
        {2'b01, 2'b10, 5'd28}     : data <= {5'd10, 5'd5};
        {2'b01, 2'b10, 5'd29}     : data <= {5'd11, 5'd3};
        {2'b01, 2'b10, 5'd30}     : data <= {5'd11, 5'd1};
        {2'b01, 2'b10, 5'd31}     : data <= {5'd11, -5'd1};
        
        {2'b01, 2'b00, 5'd0}      : data <= {5'd11, 5'd4};
        {2'b01, 2'b00, 5'd1}      : data <= {5'd11, 5'd1};
        {2'b01, 2'b00, 5'd2}      : data <= {5'd11, -5'd1};
        {2'b01, 2'b00, 5'd3}      : data <= {5'd11, -5'd3};
        {2'b01, 2'b00, 5'd4}      : data <= {5'd10, -5'd5};
        {2'b01, 2'b00, 5'd5}      : data <= {5'd9, -5'd7};
        {2'b01, 2'b00, 5'd6}      : data <= {5'd7, -5'd8};
        {2'b01, 2'b00, 5'd7}      : data <= {5'd6, -5'd10};
        {2'b01, 2'b00, 5'd8}      : data <= {5'd4, -5'd11};
        {2'b01, 2'b00, 5'd9}      : data <= {5'd1, -5'd11};
        {2'b01, 2'b00, 5'd10}     : data <= {-5'd1, -5'd11};
        {2'b01, 2'b00, 5'd11}     : data <= {-5'd3, -5'd11};
        {2'b01, 2'b00, 5'd12}     : data <= {-5'd5, -5'd10};
        {2'b01, 2'b00, 5'd13}     : data <= {-5'd7, -5'd9};
        {2'b01, 2'b00, 5'd14}     : data <= {-5'd8, -5'd7};
        {2'b01, 2'b00, 5'd15}     : data <= {-5'd10, -5'd6};
        {2'b01, 2'b00, 5'd16}     : data <= {-5'd11, -5'd4};
        {2'b01, 2'b00, 5'd17}     : data <= {-5'd11, -5'd1};
        {2'b01, 2'b00, 5'd18}     : data <= {-5'd11, 5'd1};
        {2'b01, 2'b00, 5'd19}     : data <= {-5'd11, 5'd3};
        {2'b01, 2'b00, 5'd20}     : data <= {-5'd10, 5'd5};
        {2'b01, 2'b00, 5'd21}     : data <= {-5'd9, 5'd7};
        {2'b01, 2'b00, 5'd22}     : data <= {-5'd7, 5'd8};
        {2'b01, 2'b00, 5'd23}     : data <= {-5'd6, 5'd10};
        {2'b01, 2'b00, 5'd24}     : data <= {-5'd4, 5'd11};
        {2'b01, 2'b00, 5'd25}     : data <= {-5'd1, 5'd11};
        {2'b01, 2'b00, 5'd26}     : data <= {5'd1, 5'd11};
        {2'b01, 2'b00, 5'd27}     : data <= {5'd3, 5'd11};
        {2'b01, 2'b00, 5'd28}     : data <= {5'd5, 5'd10};
        {2'b01, 2'b00, 5'd29}     : data <= {5'd7, 5'd9};
        {2'b01, 2'b00, 5'd30}     : data <= {5'd8, 5'd7};
        {2'b01, 2'b00, 5'd31}     : data <= {5'd10, 5'd6};
        
        {2'b01, 2'b01, 5'd0}      : data <= {5'd11, 5'd11};
        {2'b01, 2'b01, 5'd1}      : data <= {5'd12, 5'd8};
        {2'b01, 2'b01, 5'd2}      : data <= {5'd14, 5'd6};
        {2'b01, 2'b01, 5'd3}      : data <= {5'd15, 5'd3};
        {2'b01, 2'b01, 5'd4}      : data <= {5'd15, 5'd0};
        {2'b01, 2'b01, 5'd5}      : data <= {5'd15, -5'd3};
        {2'b01, 2'b01, 5'd6}      : data <= {5'd14, -5'd6};
        {2'b01, 2'b01, 5'd7}      : data <= {5'd12, -5'd8};
        {2'b01, 2'b01, 5'd8}      : data <= {5'd11, -5'd11};
        {2'b01, 2'b01, 5'd9}      : data <= {5'd8, -5'd12};
        {2'b01, 2'b01, 5'd10}     : data <= {5'd6, -5'd14};
        {2'b01, 2'b01, 5'd11}     : data <= {5'd3, -5'd15};
        {2'b01, 2'b01, 5'd12}     : data <= {5'd0, -5'd15};
        {2'b01, 2'b01, 5'd13}     : data <= {-5'd3, -5'd15};
        {2'b01, 2'b01, 5'd14}     : data <= {-5'd6, -5'd14};
        {2'b01, 2'b01, 5'd15}     : data <= {-5'd8, -5'd12};
        {2'b01, 2'b01, 5'd16}     : data <= {-5'd11, -5'd11};
        {2'b01, 2'b01, 5'd17}     : data <= {-5'd12, -5'd8};
        {2'b01, 2'b01, 5'd18}     : data <= {-5'd14, -5'd6};
        {2'b01, 2'b01, 5'd19}     : data <= {-5'd15, -5'd3};
        {2'b01, 2'b01, 5'd20}     : data <= {-5'd15, 5'd0};
        {2'b01, 2'b01, 5'd21}     : data <= {-5'd15, 5'd3};
        {2'b01, 2'b01, 5'd22}     : data <= {-5'd14, 5'd6};
        {2'b01, 2'b01, 5'd23}     : data <= {-5'd12, 5'd8};
        {2'b01, 2'b01, 5'd24}     : data <= {-5'd11, 5'd11};
        {2'b01, 2'b01, 5'd25}     : data <= {-5'd8, 5'd12};
        {2'b01, 2'b01, 5'd26}     : data <= {-5'd6, 5'd14};
        {2'b01, 2'b01, 5'd27}     : data <= {-5'd3, 5'd15};
        {2'b01, 2'b01, 5'd28}     : data <= {5'd0, 5'd15};
        {2'b01, 2'b01, 5'd29}     : data <= {5'd3, 5'd15};
        {2'b01, 2'b01, 5'd30}     : data <= {5'd6, 5'd14};
        {2'b01, 2'b01, 5'd31}     : data <= {5'd8, 5'd12};
    endcase
end

endmodule