`ifndef ID_DB_SVH
`define ID_DB_SVH

struct {
    int  acq_freq_shift;
    int  acq_prestore;
    int  max_args;
    int  dds_sin_cos;
    int  dds_bin;
    int  acq_bram_controller;
    int  fsm_acq_controller;
    int  acq_ip;
    int  connectbus;
    int  time_ch;
    int  axi_trig;
    int  z706_deser;
    int  psp_gen;
    int  irq_ctrl;
    int  corr_ch;
    int  oryx;
    int  sigmag_test;
    int  bdss;
    int  data_collector;
    int  trcv;
    int  time_com;
    int  ref_in_interpretator;
    int  calibration;
    int  stuff;
    int  frequency_counter;
    int  RGB;
    int  cmpo_deser;
    int  axi_performance;
    int  axi_hp_performance;
    int  axi_hp_master;
    int  cov_matrix;
    int  crpa_old;
    int  null_former;
    int  crpa;
    int  XADC_7000;
    int  imi_channel;
    int  vitterby_dec;
    int  gps_ca_prn_gen;
    int  FIR;
    int  HETERODYNE;
    int  cvm_ram;
    int  imitator;
    int  dma_intbus_axi_hp;
    int  empty;
    int  axi_uartlite_spi;
    int  axi_uart;
    int  data_recorder;
    int  adc_interconnect;
    int  decimator;
    int  samtec_ddr_decoder;
    int  cspp_adc_deser;
    int  cspp;
    int  prn_ram;
    int  dma;
    int  mem_controller;
    int  fir_syst;
    int  prn_gen_facq;
    int  facq_prn_ram;
    int  dsp_lut_iq;
    int  normalizer;
    int  acq_fft_IP;
    int  prn_gen_facq_fft;
    int  prestore_fft;
    int  lim_cntr;
    int  heterodyne_up;
} ID_DB = '{
    16'h19BE,// acq_freq_shift
    16'hAB2C,// acq_prestore
    16'h1760,// max_args
    16'h6237,// dds_sin_cos
    16'h4E46,// dds_bin
    16'h655C,// acq_bram_controller
    16'hF646,// fsm_acq_controller
    16'h18F8,// acq_ip
    16'h46E4,// connectbus
    16'h74,// time_ch
    16'hD090,// axi_trig
    16'hE7E1,// z706_deser
    16'h37,// psp_gen
    16'h11,// irq_ctrl
    16'hAB13,// corr_ch
    16'hD8DC,// oryx
    16'hE004,// sigmag_test
    16'h2082,// bdss
    16'hB0BA,// data_collector
    16'hD627,// trcv
    16'hE9D2,// time_com
    16'hA1E1,// ref_in_interpretator
    16'h474B,// calibration
    16'h1FE9,// stuff
    16'h1C40,// frequency_counter
    16'h8BFF,// RGB
    16'hB1AA,// cmpo_deser
    16'hF51E,// axi_performance
    16'hF701,// axi_hp_performance
    16'h2859,// axi_hp_master
    16'hF877,// cov_matrix
    16'hF507,// crpa_old
    16'h7C41,// null_former
    16'hCCDE,// crpa
    16'h2452,// XADC_7000
    16'h6BF8,// imi_channel
    16'hEA6C,// vitterby_dec
    16'hCACD,// gps_ca_prn_gen
    16'hF5A0,// FIR
    16'hA7DD,// HETERODYNE
    16'h924,// cvm_ram
    16'hD95F,// imitator
    16'hEF19,// dma_intbus_axi_hp
    16'h0,// empty
    16'hADC0,// axi_uartlite_spi
    16'hC1FA,// axi_uart
    16'hB0BE,// data_recorder
    16'hBE3D,// adc_interconnect
    16'h6468,// decimator
    16'hA7CC,// samtec_ddr_decoder
    16'h2BD2,// cspp_adc_deser
    16'hB4BE,// cspp
    16'h826,// prn_ram
    16'hBD1,// dma
    16'h6756,// mem_controller
    16'h18DD,// fir_syst
    16'hD2CD,// prn_gen_facq
    16'hCE4E,// facq_prn_ram
    16'hB1DF,// dsp_lut_iq
    16'h512D,// normalizer
    16'hF6EB,// acq_fft_IP
    16'hAA8F,// prn_gen_facq_fft
    16'hB9E4,// prestore_fft
    16'hF340,// lim_cntr
    16'h8D1 // heterodyne_up
};

`endif
